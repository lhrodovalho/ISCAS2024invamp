magic
tech gf180mcuC
timestamp 1697147137
<< nwell >>
rect -24 270 1068 474
<< nmos >>
rect 0 12 12 48
rect 24 12 36 48
rect 48 12 60 48
rect 72 12 84 48
rect 96 12 108 48
rect 120 12 132 48
rect 144 12 156 48
rect 168 12 180 48
rect 216 12 228 48
rect 240 12 252 48
rect 264 12 276 48
rect 288 12 300 48
rect 312 12 324 48
rect 336 12 348 48
rect 360 12 372 48
rect 384 12 396 48
rect 432 12 444 48
rect 456 12 468 48
rect 480 12 492 48
rect 504 12 516 48
rect 528 12 540 48
rect 552 12 564 48
rect 576 12 588 48
rect 600 12 612 48
rect 648 12 660 48
rect 672 12 684 48
rect 696 12 708 48
rect 720 12 732 48
rect 744 12 756 48
rect 768 12 780 48
rect 792 12 804 48
rect 816 12 828 48
rect 864 12 876 48
rect 888 12 900 48
rect 912 12 924 48
rect 936 12 948 48
rect 960 12 972 48
rect 984 12 996 48
rect 1008 12 1020 48
rect 1032 12 1044 48
rect 1080 12 1092 48
rect 1104 12 1116 48
rect 1128 12 1140 48
rect 1152 12 1164 48
rect 1176 12 1188 48
rect 1200 12 1212 48
rect 1224 12 1236 48
rect 1248 12 1260 48
<< mvnmos >>
rect 0 180 12 216
rect 24 180 36 216
rect 48 180 60 216
rect 72 180 84 216
rect 96 180 108 216
rect 120 180 132 216
rect 144 180 156 216
rect 168 180 180 216
rect 216 180 228 216
rect 240 180 252 216
rect 264 180 276 216
rect 288 180 300 216
rect 312 180 324 216
rect 336 180 348 216
rect 360 180 372 216
rect 384 180 396 216
rect 432 180 444 216
rect 456 180 468 216
rect 480 180 492 216
rect 504 180 516 216
rect 528 180 540 216
rect 552 180 564 216
rect 576 180 588 216
rect 600 180 612 216
rect 648 180 660 216
rect 672 180 684 216
rect 696 180 708 216
rect 720 180 732 216
rect 744 180 756 216
rect 768 180 780 216
rect 792 180 804 216
rect 816 180 828 216
rect 864 180 876 216
rect 912 180 924 216
rect 936 180 948 216
rect 960 180 972 216
rect 984 180 996 216
rect 1008 180 1020 216
rect 1032 180 1044 216
rect 1080 180 1092 216
rect 1104 180 1116 216
rect 1128 180 1140 216
rect 1152 180 1164 216
rect 1176 180 1188 216
rect 1200 180 1212 216
rect 1224 180 1236 216
rect 1248 180 1260 216
<< mvpmos >>
rect 0 408 12 444
rect 24 408 36 444
rect 48 408 60 444
rect 72 408 84 444
rect 96 408 108 444
rect 120 408 132 444
rect 144 408 156 444
rect 168 408 180 444
rect 216 408 228 444
rect 240 408 252 444
rect 264 408 276 444
rect 288 408 300 444
rect 312 408 324 444
rect 336 408 348 444
rect 360 408 372 444
rect 384 408 396 444
rect 432 408 444 444
rect 456 408 468 444
rect 480 408 492 444
rect 504 408 516 444
rect 528 408 540 444
rect 552 408 564 444
rect 576 408 588 444
rect 600 408 612 444
rect 648 408 660 444
rect 672 408 684 444
rect 696 408 708 444
rect 720 408 732 444
rect 744 408 756 444
rect 768 408 780 444
rect 792 408 804 444
rect 816 408 828 444
rect 864 408 876 444
rect 888 408 900 444
rect 912 408 924 444
rect 936 408 948 444
rect 960 408 972 444
rect 984 408 996 444
rect 1008 408 1020 444
rect 1032 408 1044 444
rect 0 324 12 360
rect 24 324 36 360
rect 48 324 60 360
rect 72 324 84 360
rect 96 324 108 360
rect 120 324 132 360
rect 144 324 156 360
rect 168 324 180 360
rect 216 324 228 360
rect 240 324 252 360
rect 264 324 276 360
rect 288 324 300 360
rect 312 324 324 360
rect 336 324 348 360
rect 360 324 372 360
rect 384 324 396 360
rect 432 324 444 360
rect 456 324 468 360
rect 480 324 492 360
rect 504 324 516 360
rect 528 324 540 360
rect 552 324 564 360
rect 576 324 588 360
rect 600 324 612 360
rect 648 324 660 360
rect 672 324 684 360
rect 696 324 708 360
rect 720 324 732 360
rect 744 324 756 360
rect 768 324 780 360
rect 792 324 804 360
rect 816 324 828 360
rect 864 324 876 360
rect 888 324 900 360
rect 912 324 924 360
rect 936 324 948 360
rect 960 324 972 360
rect 984 324 996 360
rect 1008 324 1020 360
rect 1032 324 1044 360
<< ndiff >>
rect -12 45 0 48
rect -12 39 -9 45
rect -3 39 0 45
rect -12 33 0 39
rect -12 27 -9 33
rect -3 27 0 33
rect -12 21 0 27
rect -12 15 -9 21
rect -3 15 0 21
rect -12 12 0 15
rect 12 12 24 48
rect 36 45 48 48
rect 36 39 39 45
rect 45 39 48 45
rect 36 33 48 39
rect 36 27 39 33
rect 45 27 48 33
rect 36 21 48 27
rect 36 15 39 21
rect 45 15 48 21
rect 36 12 48 15
rect 60 12 72 48
rect 84 45 96 48
rect 84 39 87 45
rect 93 39 96 45
rect 84 33 96 39
rect 84 27 87 33
rect 93 27 96 33
rect 84 21 96 27
rect 84 15 87 21
rect 93 15 96 21
rect 84 12 96 15
rect 108 12 120 48
rect 132 45 144 48
rect 132 39 135 45
rect 141 39 144 45
rect 132 33 144 39
rect 132 27 135 33
rect 141 27 144 33
rect 132 21 144 27
rect 132 15 135 21
rect 141 15 144 21
rect 132 12 144 15
rect 156 12 168 48
rect 180 45 192 48
rect 180 39 183 45
rect 189 39 192 45
rect 180 33 192 39
rect 180 27 183 33
rect 189 27 192 33
rect 180 21 192 27
rect 180 15 183 21
rect 189 15 192 21
rect 180 12 192 15
rect 204 45 216 48
rect 204 39 207 45
rect 213 39 216 45
rect 204 33 216 39
rect 204 27 207 33
rect 213 27 216 33
rect 204 21 216 27
rect 204 15 207 21
rect 213 15 216 21
rect 204 12 216 15
rect 228 12 240 48
rect 252 45 264 48
rect 252 39 255 45
rect 261 39 264 45
rect 252 33 264 39
rect 252 27 255 33
rect 261 27 264 33
rect 252 21 264 27
rect 252 15 255 21
rect 261 15 264 21
rect 252 12 264 15
rect 276 12 288 48
rect 300 45 312 48
rect 300 39 303 45
rect 309 39 312 45
rect 300 33 312 39
rect 300 27 303 33
rect 309 27 312 33
rect 300 21 312 27
rect 300 15 303 21
rect 309 15 312 21
rect 300 12 312 15
rect 324 12 336 48
rect 348 45 360 48
rect 348 39 351 45
rect 357 39 360 45
rect 348 33 360 39
rect 348 27 351 33
rect 357 27 360 33
rect 348 21 360 27
rect 348 15 351 21
rect 357 15 360 21
rect 348 12 360 15
rect 372 12 384 48
rect 396 45 408 48
rect 396 39 399 45
rect 405 39 408 45
rect 396 33 408 39
rect 396 27 399 33
rect 405 27 408 33
rect 396 21 408 27
rect 396 15 399 21
rect 405 15 408 21
rect 396 12 408 15
rect 420 45 432 48
rect 420 39 423 45
rect 429 39 432 45
rect 420 33 432 39
rect 420 27 423 33
rect 429 27 432 33
rect 420 21 432 27
rect 420 15 423 21
rect 429 15 432 21
rect 420 12 432 15
rect 444 12 456 48
rect 468 12 480 48
rect 492 12 504 48
rect 516 45 528 48
rect 516 39 519 45
rect 525 39 528 45
rect 516 33 528 39
rect 516 27 519 33
rect 525 27 528 33
rect 516 21 528 27
rect 516 15 519 21
rect 525 15 528 21
rect 516 12 528 15
rect 540 12 552 48
rect 564 12 576 48
rect 588 12 600 48
rect 612 45 624 48
rect 612 39 615 45
rect 621 39 624 45
rect 612 33 624 39
rect 612 27 615 33
rect 621 27 624 33
rect 612 21 624 27
rect 612 15 615 21
rect 621 15 624 21
rect 612 12 624 15
rect 636 45 648 48
rect 636 39 639 45
rect 645 39 648 45
rect 636 33 648 39
rect 636 27 639 33
rect 645 27 648 33
rect 636 21 648 27
rect 636 15 639 21
rect 645 15 648 21
rect 636 12 648 15
rect 660 12 672 48
rect 684 12 696 48
rect 708 12 720 48
rect 732 45 744 48
rect 732 39 735 45
rect 741 39 744 45
rect 732 33 744 39
rect 732 27 735 33
rect 741 27 744 33
rect 732 21 744 27
rect 732 15 735 21
rect 741 15 744 21
rect 732 12 744 15
rect 756 12 768 48
rect 780 12 792 48
rect 804 12 816 48
rect 828 45 840 48
rect 828 39 831 45
rect 837 39 840 45
rect 828 33 840 39
rect 828 27 831 33
rect 837 27 840 33
rect 828 21 840 27
rect 828 15 831 21
rect 837 15 840 21
rect 828 12 840 15
rect 852 45 864 48
rect 852 39 855 45
rect 861 39 864 45
rect 852 33 864 39
rect 852 27 855 33
rect 861 27 864 33
rect 852 21 864 27
rect 852 15 855 21
rect 861 15 864 21
rect 852 12 864 15
rect 876 12 888 48
rect 900 12 912 48
rect 924 12 936 48
rect 948 12 960 48
rect 972 12 984 48
rect 996 12 1008 48
rect 1020 12 1032 48
rect 1044 45 1056 48
rect 1044 39 1047 45
rect 1053 39 1056 45
rect 1044 33 1056 39
rect 1044 27 1047 33
rect 1053 27 1056 33
rect 1044 21 1056 27
rect 1044 15 1047 21
rect 1053 15 1056 21
rect 1044 12 1056 15
rect 1068 45 1080 48
rect 1068 39 1071 45
rect 1077 39 1080 45
rect 1068 33 1080 39
rect 1068 27 1071 33
rect 1077 27 1080 33
rect 1068 21 1080 27
rect 1068 15 1071 21
rect 1077 15 1080 21
rect 1068 12 1080 15
rect 1092 12 1104 48
rect 1116 12 1128 48
rect 1140 12 1152 48
rect 1164 45 1176 48
rect 1164 39 1167 45
rect 1173 39 1176 45
rect 1164 33 1176 39
rect 1164 27 1167 33
rect 1173 27 1176 33
rect 1164 21 1176 27
rect 1164 15 1167 21
rect 1173 15 1176 21
rect 1164 12 1176 15
rect 1188 12 1200 48
rect 1212 12 1224 48
rect 1236 12 1248 48
rect 1260 45 1272 48
rect 1260 39 1263 45
rect 1269 39 1272 45
rect 1260 33 1272 39
rect 1260 27 1263 33
rect 1269 27 1272 33
rect 1260 21 1272 27
rect 1260 15 1263 21
rect 1269 15 1272 21
rect 1260 12 1272 15
<< mvndiff >>
rect -12 213 0 216
rect -12 207 -9 213
rect -3 207 0 213
rect -12 201 0 207
rect -12 195 -9 201
rect -3 195 0 201
rect -12 189 0 195
rect -12 183 -9 189
rect -3 183 0 189
rect -12 180 0 183
rect 12 213 24 216
rect 12 207 15 213
rect 21 207 24 213
rect 12 201 24 207
rect 12 195 15 201
rect 21 195 24 201
rect 12 189 24 195
rect 12 183 15 189
rect 21 183 24 189
rect 12 180 24 183
rect 36 213 48 216
rect 36 207 39 213
rect 45 207 48 213
rect 36 201 48 207
rect 36 195 39 201
rect 45 195 48 201
rect 36 189 48 195
rect 36 183 39 189
rect 45 183 48 189
rect 36 180 48 183
rect 60 213 72 216
rect 60 207 63 213
rect 69 207 72 213
rect 60 201 72 207
rect 60 195 63 201
rect 69 195 72 201
rect 60 189 72 195
rect 60 183 63 189
rect 69 183 72 189
rect 60 180 72 183
rect 84 213 96 216
rect 84 207 87 213
rect 93 207 96 213
rect 84 201 96 207
rect 84 195 87 201
rect 93 195 96 201
rect 84 189 96 195
rect 84 183 87 189
rect 93 183 96 189
rect 84 180 96 183
rect 108 213 120 216
rect 108 207 111 213
rect 117 207 120 213
rect 108 201 120 207
rect 108 195 111 201
rect 117 195 120 201
rect 108 189 120 195
rect 108 183 111 189
rect 117 183 120 189
rect 108 180 120 183
rect 132 213 144 216
rect 132 207 135 213
rect 141 207 144 213
rect 132 201 144 207
rect 132 195 135 201
rect 141 195 144 201
rect 132 189 144 195
rect 132 183 135 189
rect 141 183 144 189
rect 132 180 144 183
rect 156 213 168 216
rect 156 207 159 213
rect 165 207 168 213
rect 156 201 168 207
rect 156 195 159 201
rect 165 195 168 201
rect 156 189 168 195
rect 156 183 159 189
rect 165 183 168 189
rect 156 180 168 183
rect 180 213 192 216
rect 180 207 183 213
rect 189 207 192 213
rect 180 201 192 207
rect 180 195 183 201
rect 189 195 192 201
rect 180 189 192 195
rect 180 183 183 189
rect 189 183 192 189
rect 180 180 192 183
rect 204 213 216 216
rect 204 207 207 213
rect 213 207 216 213
rect 204 201 216 207
rect 204 195 207 201
rect 213 195 216 201
rect 204 189 216 195
rect 204 183 207 189
rect 213 183 216 189
rect 204 180 216 183
rect 228 180 240 216
rect 252 180 264 216
rect 276 180 288 216
rect 300 213 312 216
rect 300 207 303 213
rect 309 207 312 213
rect 300 201 312 207
rect 300 195 303 201
rect 309 195 312 201
rect 300 189 312 195
rect 300 183 303 189
rect 309 183 312 189
rect 300 180 312 183
rect 324 180 336 216
rect 348 180 360 216
rect 372 180 384 216
rect 396 213 408 216
rect 396 207 399 213
rect 405 207 408 213
rect 396 201 408 207
rect 396 195 399 201
rect 405 195 408 201
rect 396 189 408 195
rect 396 183 399 189
rect 405 183 408 189
rect 396 180 408 183
rect 420 213 432 216
rect 420 207 423 213
rect 429 207 432 213
rect 420 201 432 207
rect 420 195 423 201
rect 429 195 432 201
rect 420 189 432 195
rect 420 183 423 189
rect 429 183 432 189
rect 420 180 432 183
rect 444 180 456 216
rect 468 180 480 216
rect 492 180 504 216
rect 516 213 528 216
rect 516 207 519 213
rect 525 207 528 213
rect 516 201 528 207
rect 516 195 519 201
rect 525 195 528 201
rect 516 189 528 195
rect 516 183 519 189
rect 525 183 528 189
rect 516 180 528 183
rect 540 180 552 216
rect 564 180 576 216
rect 588 180 600 216
rect 612 213 624 216
rect 612 207 615 213
rect 621 207 624 213
rect 612 201 624 207
rect 612 195 615 201
rect 621 195 624 201
rect 612 189 624 195
rect 612 183 615 189
rect 621 183 624 189
rect 612 180 624 183
rect 636 213 648 216
rect 636 207 639 213
rect 645 207 648 213
rect 636 201 648 207
rect 636 195 639 201
rect 645 195 648 201
rect 636 189 648 195
rect 636 183 639 189
rect 645 183 648 189
rect 636 180 648 183
rect 660 180 672 216
rect 684 180 696 216
rect 708 180 720 216
rect 732 213 744 216
rect 732 207 735 213
rect 741 207 744 213
rect 732 201 744 207
rect 732 195 735 201
rect 741 195 744 201
rect 732 189 744 195
rect 732 183 735 189
rect 741 183 744 189
rect 732 180 744 183
rect 756 180 768 216
rect 780 180 792 216
rect 804 180 816 216
rect 828 213 840 216
rect 828 207 831 213
rect 837 207 840 213
rect 828 201 840 207
rect 828 195 831 201
rect 837 195 840 201
rect 828 189 840 195
rect 828 183 831 189
rect 837 183 840 189
rect 828 180 840 183
rect 852 213 864 216
rect 852 207 855 213
rect 861 207 864 213
rect 852 201 864 207
rect 852 195 855 201
rect 861 195 864 201
rect 852 189 864 195
rect 852 183 855 189
rect 861 183 864 189
rect 852 180 864 183
rect 876 213 888 216
rect 876 207 879 213
rect 885 207 888 213
rect 876 201 888 207
rect 876 195 879 201
rect 885 195 888 201
rect 876 189 888 195
rect 876 183 879 189
rect 885 183 888 189
rect 876 180 888 183
rect 900 213 912 216
rect 900 207 903 213
rect 909 207 912 213
rect 900 201 912 207
rect 900 195 903 201
rect 909 195 912 201
rect 900 189 912 195
rect 900 183 903 189
rect 909 183 912 189
rect 900 180 912 183
rect 924 180 936 216
rect 948 180 960 216
rect 972 180 984 216
rect 996 180 1008 216
rect 1020 180 1032 216
rect 1044 213 1056 216
rect 1044 207 1047 213
rect 1053 207 1056 213
rect 1044 201 1056 207
rect 1044 195 1047 201
rect 1053 195 1056 201
rect 1044 189 1056 195
rect 1044 183 1047 189
rect 1053 183 1056 189
rect 1044 180 1056 183
rect 1068 213 1080 216
rect 1068 207 1071 213
rect 1077 207 1080 213
rect 1068 201 1080 207
rect 1068 195 1071 201
rect 1077 195 1080 201
rect 1068 189 1080 195
rect 1068 183 1071 189
rect 1077 183 1080 189
rect 1068 180 1080 183
rect 1092 180 1104 216
rect 1116 180 1128 216
rect 1140 180 1152 216
rect 1164 213 1176 216
rect 1164 207 1167 213
rect 1173 207 1176 213
rect 1164 201 1176 207
rect 1164 195 1167 201
rect 1173 195 1176 201
rect 1164 189 1176 195
rect 1164 183 1167 189
rect 1173 183 1176 189
rect 1164 180 1176 183
rect 1188 180 1200 216
rect 1212 180 1224 216
rect 1236 180 1248 216
rect 1260 213 1272 216
rect 1260 207 1263 213
rect 1269 207 1272 213
rect 1260 201 1272 207
rect 1260 195 1263 201
rect 1269 195 1272 201
rect 1260 189 1272 195
rect 1260 183 1263 189
rect 1269 183 1272 189
rect 1260 180 1272 183
<< mvpdiff >>
rect -12 441 0 444
rect -12 435 -9 441
rect -3 435 0 441
rect -12 429 0 435
rect -12 423 -9 429
rect -3 423 0 429
rect -12 417 0 423
rect -12 411 -9 417
rect -3 411 0 417
rect -12 408 0 411
rect 12 441 24 444
rect 12 435 15 441
rect 21 435 24 441
rect 12 429 24 435
rect 12 423 15 429
rect 21 423 24 429
rect 12 417 24 423
rect 12 411 15 417
rect 21 411 24 417
rect 12 408 24 411
rect 36 441 48 444
rect 36 435 39 441
rect 45 435 48 441
rect 36 429 48 435
rect 36 423 39 429
rect 45 423 48 429
rect 36 417 48 423
rect 36 411 39 417
rect 45 411 48 417
rect 36 408 48 411
rect 60 441 72 444
rect 60 435 63 441
rect 69 435 72 441
rect 60 429 72 435
rect 60 423 63 429
rect 69 423 72 429
rect 60 417 72 423
rect 60 411 63 417
rect 69 411 72 417
rect 60 408 72 411
rect 84 441 96 444
rect 84 435 87 441
rect 93 435 96 441
rect 84 429 96 435
rect 84 423 87 429
rect 93 423 96 429
rect 84 417 96 423
rect 84 411 87 417
rect 93 411 96 417
rect 84 408 96 411
rect 108 441 120 444
rect 108 435 111 441
rect 117 435 120 441
rect 108 429 120 435
rect 108 423 111 429
rect 117 423 120 429
rect 108 417 120 423
rect 108 411 111 417
rect 117 411 120 417
rect 108 408 120 411
rect 132 441 144 444
rect 132 435 135 441
rect 141 435 144 441
rect 132 429 144 435
rect 132 423 135 429
rect 141 423 144 429
rect 132 417 144 423
rect 132 411 135 417
rect 141 411 144 417
rect 132 408 144 411
rect 156 441 168 444
rect 156 435 159 441
rect 165 435 168 441
rect 156 429 168 435
rect 156 423 159 429
rect 165 423 168 429
rect 156 417 168 423
rect 156 411 159 417
rect 165 411 168 417
rect 156 408 168 411
rect 180 441 192 444
rect 180 435 183 441
rect 189 435 192 441
rect 180 429 192 435
rect 180 423 183 429
rect 189 423 192 429
rect 180 417 192 423
rect 180 411 183 417
rect 189 411 192 417
rect 180 408 192 411
rect 204 441 216 444
rect 204 435 207 441
rect 213 435 216 441
rect 204 429 216 435
rect 204 423 207 429
rect 213 423 216 429
rect 204 417 216 423
rect 204 411 207 417
rect 213 411 216 417
rect 204 408 216 411
rect 228 408 240 444
rect 252 441 264 444
rect 252 435 255 441
rect 261 435 264 441
rect 252 429 264 435
rect 252 423 255 429
rect 261 423 264 429
rect 252 417 264 423
rect 252 411 255 417
rect 261 411 264 417
rect 252 408 264 411
rect 276 408 288 444
rect 300 441 312 444
rect 300 435 303 441
rect 309 435 312 441
rect 300 429 312 435
rect 300 423 303 429
rect 309 423 312 429
rect 300 417 312 423
rect 300 411 303 417
rect 309 411 312 417
rect 300 408 312 411
rect 324 408 336 444
rect 348 441 360 444
rect 348 435 351 441
rect 357 435 360 441
rect 348 429 360 435
rect 348 423 351 429
rect 357 423 360 429
rect 348 417 360 423
rect 348 411 351 417
rect 357 411 360 417
rect 348 408 360 411
rect 372 408 384 444
rect 396 441 408 444
rect 396 435 399 441
rect 405 435 408 441
rect 396 429 408 435
rect 396 423 399 429
rect 405 423 408 429
rect 396 417 408 423
rect 396 411 399 417
rect 405 411 408 417
rect 396 408 408 411
rect 420 441 432 444
rect 420 435 423 441
rect 429 435 432 441
rect 420 429 432 435
rect 420 423 423 429
rect 429 423 432 429
rect 420 417 432 423
rect 420 411 423 417
rect 429 411 432 417
rect 420 408 432 411
rect 444 408 456 444
rect 468 441 480 444
rect 468 435 471 441
rect 477 435 480 441
rect 468 429 480 435
rect 468 423 471 429
rect 477 423 480 429
rect 468 417 480 423
rect 468 411 471 417
rect 477 411 480 417
rect 468 408 480 411
rect 492 408 504 444
rect 516 441 528 444
rect 516 435 519 441
rect 525 435 528 441
rect 516 429 528 435
rect 516 423 519 429
rect 525 423 528 429
rect 516 417 528 423
rect 516 411 519 417
rect 525 411 528 417
rect 516 408 528 411
rect 540 408 552 444
rect 564 441 576 444
rect 564 435 567 441
rect 573 435 576 441
rect 564 429 576 435
rect 564 423 567 429
rect 573 423 576 429
rect 564 417 576 423
rect 564 411 567 417
rect 573 411 576 417
rect 564 408 576 411
rect 588 408 600 444
rect 612 441 624 444
rect 612 435 615 441
rect 621 435 624 441
rect 612 429 624 435
rect 612 423 615 429
rect 621 423 624 429
rect 612 417 624 423
rect 612 411 615 417
rect 621 411 624 417
rect 612 408 624 411
rect 636 441 648 444
rect 636 435 639 441
rect 645 435 648 441
rect 636 429 648 435
rect 636 423 639 429
rect 645 423 648 429
rect 636 417 648 423
rect 636 411 639 417
rect 645 411 648 417
rect 636 408 648 411
rect 660 408 672 444
rect 684 408 696 444
rect 708 408 720 444
rect 732 408 744 444
rect 756 408 768 444
rect 780 408 792 444
rect 804 408 816 444
rect 828 441 840 444
rect 828 435 831 441
rect 837 435 840 441
rect 828 429 840 435
rect 828 423 831 429
rect 837 423 840 429
rect 828 417 840 423
rect 828 411 831 417
rect 837 411 840 417
rect 828 408 840 411
rect 852 441 864 444
rect 852 435 855 441
rect 861 435 864 441
rect 852 429 864 435
rect 852 423 855 429
rect 861 423 864 429
rect 852 417 864 423
rect 852 411 855 417
rect 861 411 864 417
rect 852 408 864 411
rect 876 408 888 444
rect 900 408 912 444
rect 924 408 936 444
rect 948 408 960 444
rect 972 408 984 444
rect 996 408 1008 444
rect 1020 408 1032 444
rect 1044 441 1056 444
rect 1044 435 1047 441
rect 1053 435 1056 441
rect 1044 429 1056 435
rect 1044 423 1047 429
rect 1053 423 1056 429
rect 1044 417 1056 423
rect 1044 411 1047 417
rect 1053 411 1056 417
rect 1044 408 1056 411
rect -12 357 0 360
rect -12 351 -9 357
rect -3 351 0 357
rect -12 345 0 351
rect -12 339 -9 345
rect -3 339 0 345
rect -12 333 0 339
rect -12 327 -9 333
rect -3 327 0 333
rect -12 324 0 327
rect 12 357 24 360
rect 12 351 15 357
rect 21 351 24 357
rect 12 345 24 351
rect 12 339 15 345
rect 21 339 24 345
rect 12 333 24 339
rect 12 327 15 333
rect 21 327 24 333
rect 12 324 24 327
rect 36 357 48 360
rect 36 351 39 357
rect 45 351 48 357
rect 36 345 48 351
rect 36 339 39 345
rect 45 339 48 345
rect 36 333 48 339
rect 36 327 39 333
rect 45 327 48 333
rect 36 324 48 327
rect 60 357 72 360
rect 60 351 63 357
rect 69 351 72 357
rect 60 345 72 351
rect 60 339 63 345
rect 69 339 72 345
rect 60 333 72 339
rect 60 327 63 333
rect 69 327 72 333
rect 60 324 72 327
rect 84 357 96 360
rect 84 351 87 357
rect 93 351 96 357
rect 84 345 96 351
rect 84 339 87 345
rect 93 339 96 345
rect 84 333 96 339
rect 84 327 87 333
rect 93 327 96 333
rect 84 324 96 327
rect 108 357 120 360
rect 108 351 111 357
rect 117 351 120 357
rect 108 345 120 351
rect 108 339 111 345
rect 117 339 120 345
rect 108 333 120 339
rect 108 327 111 333
rect 117 327 120 333
rect 108 324 120 327
rect 132 357 144 360
rect 132 351 135 357
rect 141 351 144 357
rect 132 345 144 351
rect 132 339 135 345
rect 141 339 144 345
rect 132 333 144 339
rect 132 327 135 333
rect 141 327 144 333
rect 132 324 144 327
rect 156 357 168 360
rect 156 351 159 357
rect 165 351 168 357
rect 156 345 168 351
rect 156 339 159 345
rect 165 339 168 345
rect 156 333 168 339
rect 156 327 159 333
rect 165 327 168 333
rect 156 324 168 327
rect 180 357 192 360
rect 180 351 183 357
rect 189 351 192 357
rect 180 345 192 351
rect 180 339 183 345
rect 189 339 192 345
rect 180 333 192 339
rect 180 327 183 333
rect 189 327 192 333
rect 180 324 192 327
rect 204 357 216 360
rect 204 351 207 357
rect 213 351 216 357
rect 204 345 216 351
rect 204 339 207 345
rect 213 339 216 345
rect 204 333 216 339
rect 204 327 207 333
rect 213 327 216 333
rect 204 324 216 327
rect 228 324 240 360
rect 252 357 264 360
rect 252 351 255 357
rect 261 351 264 357
rect 252 345 264 351
rect 252 339 255 345
rect 261 339 264 345
rect 252 333 264 339
rect 252 327 255 333
rect 261 327 264 333
rect 252 324 264 327
rect 276 324 288 360
rect 300 357 312 360
rect 300 351 303 357
rect 309 351 312 357
rect 300 345 312 351
rect 300 339 303 345
rect 309 339 312 345
rect 300 333 312 339
rect 300 327 303 333
rect 309 327 312 333
rect 300 324 312 327
rect 324 324 336 360
rect 348 357 360 360
rect 348 351 351 357
rect 357 351 360 357
rect 348 345 360 351
rect 348 339 351 345
rect 357 339 360 345
rect 348 333 360 339
rect 348 327 351 333
rect 357 327 360 333
rect 348 324 360 327
rect 372 324 384 360
rect 396 357 408 360
rect 396 351 399 357
rect 405 351 408 357
rect 396 345 408 351
rect 396 339 399 345
rect 405 339 408 345
rect 396 333 408 339
rect 396 327 399 333
rect 405 327 408 333
rect 396 324 408 327
rect 420 357 432 360
rect 420 351 423 357
rect 429 351 432 357
rect 420 345 432 351
rect 420 339 423 345
rect 429 339 432 345
rect 420 333 432 339
rect 420 327 423 333
rect 429 327 432 333
rect 420 324 432 327
rect 444 324 456 360
rect 468 357 480 360
rect 468 351 471 357
rect 477 351 480 357
rect 468 345 480 351
rect 468 339 471 345
rect 477 339 480 345
rect 468 333 480 339
rect 468 327 471 333
rect 477 327 480 333
rect 468 324 480 327
rect 492 324 504 360
rect 516 357 528 360
rect 516 351 519 357
rect 525 351 528 357
rect 516 345 528 351
rect 516 339 519 345
rect 525 339 528 345
rect 516 333 528 339
rect 516 327 519 333
rect 525 327 528 333
rect 516 324 528 327
rect 540 324 552 360
rect 564 357 576 360
rect 564 351 567 357
rect 573 351 576 357
rect 564 345 576 351
rect 564 339 567 345
rect 573 339 576 345
rect 564 333 576 339
rect 564 327 567 333
rect 573 327 576 333
rect 564 324 576 327
rect 588 324 600 360
rect 612 357 624 360
rect 612 351 615 357
rect 621 351 624 357
rect 612 345 624 351
rect 612 339 615 345
rect 621 339 624 345
rect 612 333 624 339
rect 612 327 615 333
rect 621 327 624 333
rect 612 324 624 327
rect 636 357 648 360
rect 636 351 639 357
rect 645 351 648 357
rect 636 345 648 351
rect 636 339 639 345
rect 645 339 648 345
rect 636 333 648 339
rect 636 327 639 333
rect 645 327 648 333
rect 636 324 648 327
rect 660 324 672 360
rect 684 324 696 360
rect 708 324 720 360
rect 732 324 744 360
rect 756 324 768 360
rect 780 324 792 360
rect 804 324 816 360
rect 828 357 840 360
rect 828 351 831 357
rect 837 351 840 357
rect 828 345 840 351
rect 828 339 831 345
rect 837 339 840 345
rect 828 333 840 339
rect 828 327 831 333
rect 837 327 840 333
rect 828 324 840 327
rect 852 357 864 360
rect 852 351 855 357
rect 861 351 864 357
rect 852 345 864 351
rect 852 339 855 345
rect 861 339 864 345
rect 852 333 864 339
rect 852 327 855 333
rect 861 327 864 333
rect 852 324 864 327
rect 876 324 888 360
rect 900 324 912 360
rect 924 324 936 360
rect 948 324 960 360
rect 972 324 984 360
rect 996 324 1008 360
rect 1020 324 1032 360
rect 1044 357 1056 360
rect 1044 351 1047 357
rect 1053 351 1056 357
rect 1044 345 1056 351
rect 1044 339 1047 345
rect 1053 339 1056 345
rect 1044 333 1056 339
rect 1044 327 1047 333
rect 1053 327 1056 333
rect 1044 324 1056 327
<< ndiffc >>
rect -9 39 -3 45
rect -9 27 -3 33
rect -9 15 -3 21
rect 39 39 45 45
rect 39 27 45 33
rect 39 15 45 21
rect 87 39 93 45
rect 87 27 93 33
rect 87 15 93 21
rect 135 39 141 45
rect 135 27 141 33
rect 135 15 141 21
rect 183 39 189 45
rect 183 27 189 33
rect 183 15 189 21
rect 207 39 213 45
rect 207 27 213 33
rect 207 15 213 21
rect 255 39 261 45
rect 255 27 261 33
rect 255 15 261 21
rect 303 39 309 45
rect 303 27 309 33
rect 303 15 309 21
rect 351 39 357 45
rect 351 27 357 33
rect 351 15 357 21
rect 399 39 405 45
rect 399 27 405 33
rect 399 15 405 21
rect 423 39 429 45
rect 423 27 429 33
rect 423 15 429 21
rect 519 39 525 45
rect 519 27 525 33
rect 519 15 525 21
rect 615 39 621 45
rect 615 27 621 33
rect 615 15 621 21
rect 639 39 645 45
rect 639 27 645 33
rect 639 15 645 21
rect 735 39 741 45
rect 735 27 741 33
rect 735 15 741 21
rect 831 39 837 45
rect 831 27 837 33
rect 831 15 837 21
rect 855 39 861 45
rect 855 27 861 33
rect 855 15 861 21
rect 1047 39 1053 45
rect 1047 27 1053 33
rect 1047 15 1053 21
rect 1071 39 1077 45
rect 1071 27 1077 33
rect 1071 15 1077 21
rect 1167 39 1173 45
rect 1167 27 1173 33
rect 1167 15 1173 21
rect 1263 39 1269 45
rect 1263 27 1269 33
rect 1263 15 1269 21
<< mvndiffc >>
rect -9 207 -3 213
rect -9 195 -3 201
rect -9 183 -3 189
rect 15 207 21 213
rect 15 195 21 201
rect 15 183 21 189
rect 39 207 45 213
rect 39 195 45 201
rect 39 183 45 189
rect 63 207 69 213
rect 63 195 69 201
rect 63 183 69 189
rect 87 207 93 213
rect 87 195 93 201
rect 87 183 93 189
rect 111 207 117 213
rect 111 195 117 201
rect 111 183 117 189
rect 135 207 141 213
rect 135 195 141 201
rect 135 183 141 189
rect 159 207 165 213
rect 159 195 165 201
rect 159 183 165 189
rect 183 207 189 213
rect 183 195 189 201
rect 183 183 189 189
rect 207 207 213 213
rect 207 195 213 201
rect 207 183 213 189
rect 303 207 309 213
rect 303 195 309 201
rect 303 183 309 189
rect 399 207 405 213
rect 399 195 405 201
rect 399 183 405 189
rect 423 207 429 213
rect 423 195 429 201
rect 423 183 429 189
rect 519 207 525 213
rect 519 195 525 201
rect 519 183 525 189
rect 615 207 621 213
rect 615 195 621 201
rect 615 183 621 189
rect 639 207 645 213
rect 639 195 645 201
rect 639 183 645 189
rect 735 207 741 213
rect 735 195 741 201
rect 735 183 741 189
rect 831 207 837 213
rect 831 195 837 201
rect 831 183 837 189
rect 855 207 861 213
rect 855 195 861 201
rect 855 183 861 189
rect 879 207 885 213
rect 879 195 885 201
rect 879 183 885 189
rect 903 207 909 213
rect 903 195 909 201
rect 903 183 909 189
rect 1047 207 1053 213
rect 1047 195 1053 201
rect 1047 183 1053 189
rect 1071 207 1077 213
rect 1071 195 1077 201
rect 1071 183 1077 189
rect 1167 207 1173 213
rect 1167 195 1173 201
rect 1167 183 1173 189
rect 1263 207 1269 213
rect 1263 195 1269 201
rect 1263 183 1269 189
<< mvpdiffc >>
rect -9 435 -3 441
rect -9 423 -3 429
rect -9 411 -3 417
rect 15 435 21 441
rect 15 423 21 429
rect 15 411 21 417
rect 39 435 45 441
rect 39 423 45 429
rect 39 411 45 417
rect 63 435 69 441
rect 63 423 69 429
rect 63 411 69 417
rect 87 435 93 441
rect 87 423 93 429
rect 87 411 93 417
rect 111 435 117 441
rect 111 423 117 429
rect 111 411 117 417
rect 135 435 141 441
rect 135 423 141 429
rect 135 411 141 417
rect 159 435 165 441
rect 159 423 165 429
rect 159 411 165 417
rect 183 435 189 441
rect 183 423 189 429
rect 183 411 189 417
rect 207 435 213 441
rect 207 423 213 429
rect 207 411 213 417
rect 255 435 261 441
rect 255 423 261 429
rect 255 411 261 417
rect 303 435 309 441
rect 303 423 309 429
rect 303 411 309 417
rect 351 435 357 441
rect 351 423 357 429
rect 351 411 357 417
rect 399 435 405 441
rect 399 423 405 429
rect 399 411 405 417
rect 423 435 429 441
rect 423 423 429 429
rect 423 411 429 417
rect 471 435 477 441
rect 471 423 477 429
rect 471 411 477 417
rect 519 435 525 441
rect 519 423 525 429
rect 519 411 525 417
rect 567 435 573 441
rect 567 423 573 429
rect 567 411 573 417
rect 615 435 621 441
rect 615 423 621 429
rect 615 411 621 417
rect 639 435 645 441
rect 639 423 645 429
rect 639 411 645 417
rect 831 435 837 441
rect 831 423 837 429
rect 831 411 837 417
rect 855 435 861 441
rect 855 423 861 429
rect 855 411 861 417
rect 1047 435 1053 441
rect 1047 423 1053 429
rect 1047 411 1053 417
rect -9 351 -3 357
rect -9 339 -3 345
rect -9 327 -3 333
rect 15 351 21 357
rect 15 339 21 345
rect 15 327 21 333
rect 39 351 45 357
rect 39 339 45 345
rect 39 327 45 333
rect 63 351 69 357
rect 63 339 69 345
rect 63 327 69 333
rect 87 351 93 357
rect 87 339 93 345
rect 87 327 93 333
rect 111 351 117 357
rect 111 339 117 345
rect 111 327 117 333
rect 135 351 141 357
rect 135 339 141 345
rect 135 327 141 333
rect 159 351 165 357
rect 159 339 165 345
rect 159 327 165 333
rect 183 351 189 357
rect 183 339 189 345
rect 183 327 189 333
rect 207 351 213 357
rect 207 339 213 345
rect 207 327 213 333
rect 255 351 261 357
rect 255 339 261 345
rect 255 327 261 333
rect 303 351 309 357
rect 303 339 309 345
rect 303 327 309 333
rect 351 351 357 357
rect 351 339 357 345
rect 351 327 357 333
rect 399 351 405 357
rect 399 339 405 345
rect 399 327 405 333
rect 423 351 429 357
rect 423 339 429 345
rect 423 327 429 333
rect 471 351 477 357
rect 471 339 477 345
rect 471 327 477 333
rect 519 351 525 357
rect 519 339 525 345
rect 519 327 525 333
rect 567 351 573 357
rect 567 339 573 345
rect 567 327 573 333
rect 615 351 621 357
rect 615 339 621 345
rect 615 327 621 333
rect 639 351 645 357
rect 639 339 645 345
rect 639 327 645 333
rect 831 351 837 357
rect 831 339 837 345
rect 831 327 837 333
rect 855 351 861 357
rect 855 339 861 345
rect 855 327 861 333
rect 1047 351 1053 357
rect 1047 339 1053 345
rect 1047 327 1053 333
<< psubdiff >>
rect -24 -3 1272 0
rect -24 -9 -21 -3
rect -15 -9 -9 -3
rect -3 -9 3 -3
rect 9 -9 15 -3
rect 21 -9 27 -3
rect 33 -9 39 -3
rect 45 -9 51 -3
rect 57 -9 63 -3
rect 69 -9 75 -3
rect 81 -9 87 -3
rect 93 -9 99 -3
rect 105 -9 111 -3
rect 117 -9 123 -3
rect 129 -9 135 -3
rect 141 -9 147 -3
rect 153 -9 159 -3
rect 165 -9 171 -3
rect 177 -9 183 -3
rect 189 -9 195 -3
rect 201 -9 207 -3
rect 213 -9 219 -3
rect 225 -9 231 -3
rect 237 -9 243 -3
rect 249 -9 255 -3
rect 261 -9 267 -3
rect 273 -9 279 -3
rect 285 -9 291 -3
rect 297 -9 303 -3
rect 309 -9 315 -3
rect 321 -9 327 -3
rect 333 -9 339 -3
rect 345 -9 351 -3
rect 357 -9 363 -3
rect 369 -9 375 -3
rect 381 -9 387 -3
rect 393 -9 399 -3
rect 405 -9 411 -3
rect 417 -9 423 -3
rect 429 -9 435 -3
rect 441 -9 447 -3
rect 453 -9 459 -3
rect 465 -9 471 -3
rect 477 -9 483 -3
rect 489 -9 495 -3
rect 501 -9 507 -3
rect 513 -9 519 -3
rect 525 -9 531 -3
rect 537 -9 543 -3
rect 549 -9 555 -3
rect 561 -9 567 -3
rect 573 -9 579 -3
rect 585 -9 591 -3
rect 597 -9 603 -3
rect 609 -9 615 -3
rect 621 -9 627 -3
rect 633 -9 639 -3
rect 645 -9 651 -3
rect 657 -9 663 -3
rect 669 -9 675 -3
rect 681 -9 687 -3
rect 693 -9 699 -3
rect 705 -9 711 -3
rect 717 -9 723 -3
rect 729 -9 735 -3
rect 741 -9 747 -3
rect 753 -9 759 -3
rect 765 -9 771 -3
rect 777 -9 783 -3
rect 789 -9 795 -3
rect 801 -9 807 -3
rect 813 -9 819 -3
rect 825 -9 831 -3
rect 837 -9 843 -3
rect 849 -9 855 -3
rect 861 -9 867 -3
rect 873 -9 879 -3
rect 885 -9 891 -3
rect 897 -9 903 -3
rect 909 -9 915 -3
rect 921 -9 927 -3
rect 933 -9 939 -3
rect 945 -9 951 -3
rect 957 -9 963 -3
rect 969 -9 975 -3
rect 981 -9 987 -3
rect 993 -9 999 -3
rect 1005 -9 1011 -3
rect 1017 -9 1023 -3
rect 1029 -9 1035 -3
rect 1041 -9 1047 -3
rect 1053 -9 1059 -3
rect 1065 -9 1071 -3
rect 1077 -9 1083 -3
rect 1089 -9 1095 -3
rect 1101 -9 1107 -3
rect 1113 -9 1119 -3
rect 1125 -9 1131 -3
rect 1137 -9 1143 -3
rect 1149 -9 1155 -3
rect 1161 -9 1167 -3
rect 1173 -9 1179 -3
rect 1185 -9 1191 -3
rect 1197 -9 1203 -3
rect 1209 -9 1215 -3
rect 1221 -9 1227 -3
rect 1233 -9 1239 -3
rect 1245 -9 1251 -3
rect 1257 -9 1263 -3
rect 1269 -9 1272 -3
rect -24 -12 1272 -9
<< mvpsubdiff >>
rect -24 261 1056 264
rect -24 255 -21 261
rect -15 255 -9 261
rect -3 255 3 261
rect 9 255 15 261
rect 21 255 27 261
rect 33 255 39 261
rect 45 255 51 261
rect 57 255 63 261
rect 69 255 75 261
rect 81 255 87 261
rect 93 255 99 261
rect 105 255 111 261
rect 117 255 123 261
rect 129 255 135 261
rect 141 255 147 261
rect 153 255 159 261
rect 165 255 171 261
rect 177 255 183 261
rect 189 255 195 261
rect 201 255 207 261
rect 213 255 219 261
rect 225 255 231 261
rect 237 255 243 261
rect 249 255 255 261
rect 261 255 267 261
rect 273 255 279 261
rect 285 255 291 261
rect 297 255 303 261
rect 309 255 315 261
rect 321 255 327 261
rect 333 255 339 261
rect 345 255 351 261
rect 357 255 363 261
rect 369 255 375 261
rect 381 255 387 261
rect 393 255 399 261
rect 405 255 411 261
rect 417 255 423 261
rect 429 255 435 261
rect 441 255 447 261
rect 453 255 459 261
rect 465 255 471 261
rect 477 255 483 261
rect 489 255 495 261
rect 501 255 507 261
rect 513 255 519 261
rect 525 255 531 261
rect 537 255 543 261
rect 549 255 555 261
rect 561 255 567 261
rect 573 255 579 261
rect 585 255 591 261
rect 597 255 603 261
rect 609 255 615 261
rect 621 255 627 261
rect 633 255 639 261
rect 645 255 651 261
rect 657 255 663 261
rect 669 255 675 261
rect 681 255 687 261
rect 693 255 699 261
rect 705 255 711 261
rect 717 255 723 261
rect 729 255 735 261
rect 741 255 747 261
rect 753 255 759 261
rect 765 255 771 261
rect 777 255 783 261
rect 789 255 795 261
rect 801 255 807 261
rect 813 255 819 261
rect 825 255 831 261
rect 837 255 843 261
rect 849 255 855 261
rect 861 255 867 261
rect 873 255 879 261
rect 885 255 891 261
rect 897 255 903 261
rect 909 255 915 261
rect 921 255 927 261
rect 933 255 939 261
rect 945 255 951 261
rect 957 255 963 261
rect 969 255 975 261
rect 981 255 987 261
rect 993 255 999 261
rect 1005 255 1011 261
rect 1017 255 1023 261
rect 1029 255 1035 261
rect 1041 255 1047 261
rect 1053 255 1056 261
rect -24 252 1056 255
<< mvnsubdiff >>
rect -12 465 1056 468
rect -12 459 -9 465
rect -3 459 3 465
rect 9 459 15 465
rect 21 459 27 465
rect 33 459 39 465
rect 45 459 51 465
rect 57 459 63 465
rect 69 459 75 465
rect 81 459 87 465
rect 93 459 99 465
rect 105 459 111 465
rect 117 459 123 465
rect 129 459 135 465
rect 141 459 147 465
rect 153 459 159 465
rect 165 459 171 465
rect 177 459 183 465
rect 189 459 195 465
rect 201 459 207 465
rect 213 459 219 465
rect 225 459 231 465
rect 237 459 243 465
rect 249 459 255 465
rect 261 459 267 465
rect 273 459 279 465
rect 285 459 291 465
rect 297 459 303 465
rect 309 459 315 465
rect 321 459 327 465
rect 333 459 339 465
rect 345 459 351 465
rect 357 459 363 465
rect 369 459 375 465
rect 381 459 387 465
rect 393 459 399 465
rect 405 459 411 465
rect 417 459 423 465
rect 429 459 435 465
rect 441 459 447 465
rect 453 459 459 465
rect 465 459 471 465
rect 477 459 483 465
rect 489 459 495 465
rect 501 459 507 465
rect 513 459 519 465
rect 525 459 531 465
rect 537 459 543 465
rect 549 459 555 465
rect 561 459 567 465
rect 573 459 579 465
rect 585 459 591 465
rect 597 459 603 465
rect 609 459 615 465
rect 621 459 627 465
rect 633 459 639 465
rect 645 459 651 465
rect 657 459 663 465
rect 669 459 675 465
rect 681 459 687 465
rect 693 459 699 465
rect 705 459 711 465
rect 717 459 723 465
rect 729 459 735 465
rect 741 459 747 465
rect 753 459 759 465
rect 765 459 771 465
rect 777 459 783 465
rect 789 459 795 465
rect 801 459 807 465
rect 813 459 819 465
rect 825 459 831 465
rect 837 459 843 465
rect 849 459 855 465
rect 861 459 867 465
rect 873 459 879 465
rect 885 459 891 465
rect 897 459 903 465
rect 909 459 915 465
rect 921 459 927 465
rect 933 459 939 465
rect 945 459 951 465
rect 957 459 963 465
rect 969 459 975 465
rect 981 459 987 465
rect 993 459 999 465
rect 1005 459 1011 465
rect 1017 459 1023 465
rect 1029 459 1035 465
rect 1041 459 1047 465
rect 1053 459 1056 465
rect -12 456 1056 459
rect -12 285 1056 288
rect -12 279 -9 285
rect -3 279 3 285
rect 9 279 15 285
rect 21 279 27 285
rect 33 279 39 285
rect 45 279 51 285
rect 57 279 63 285
rect 69 279 75 285
rect 81 279 87 285
rect 93 279 99 285
rect 105 279 111 285
rect 117 279 123 285
rect 129 279 135 285
rect 141 279 147 285
rect 153 279 159 285
rect 165 279 171 285
rect 177 279 183 285
rect 189 279 195 285
rect 201 279 207 285
rect 213 279 219 285
rect 225 279 231 285
rect 237 279 243 285
rect 249 279 255 285
rect 261 279 267 285
rect 273 279 279 285
rect 285 279 291 285
rect 297 279 303 285
rect 309 279 315 285
rect 321 279 327 285
rect 333 279 339 285
rect 345 279 351 285
rect 357 279 363 285
rect 369 279 375 285
rect 381 279 387 285
rect 393 279 399 285
rect 405 279 411 285
rect 417 279 423 285
rect 429 279 435 285
rect 441 279 447 285
rect 453 279 459 285
rect 465 279 471 285
rect 477 279 483 285
rect 489 279 495 285
rect 501 279 507 285
rect 513 279 519 285
rect 525 279 531 285
rect 537 279 543 285
rect 549 279 555 285
rect 561 279 567 285
rect 573 279 579 285
rect 585 279 591 285
rect 597 279 603 285
rect 609 279 615 285
rect 621 279 627 285
rect 633 279 639 285
rect 645 279 651 285
rect 657 279 663 285
rect 669 279 675 285
rect 681 279 687 285
rect 693 279 699 285
rect 705 279 711 285
rect 717 279 723 285
rect 729 279 735 285
rect 741 279 747 285
rect 753 279 759 285
rect 765 279 771 285
rect 777 279 783 285
rect 789 279 795 285
rect 801 279 807 285
rect 813 279 819 285
rect 825 279 831 285
rect 837 279 843 285
rect 849 279 855 285
rect 861 279 867 285
rect 873 279 879 285
rect 885 279 891 285
rect 897 279 903 285
rect 909 279 915 285
rect 921 279 927 285
rect 933 279 939 285
rect 945 279 951 285
rect 957 279 963 285
rect 969 279 975 285
rect 981 279 987 285
rect 993 279 999 285
rect 1005 279 1011 285
rect 1017 279 1023 285
rect 1029 279 1035 285
rect 1041 279 1047 285
rect 1053 279 1056 285
rect -12 276 1056 279
<< psubdiffcont >>
rect -21 -9 -15 -3
rect -9 -9 -3 -3
rect 3 -9 9 -3
rect 15 -9 21 -3
rect 27 -9 33 -3
rect 39 -9 45 -3
rect 51 -9 57 -3
rect 63 -9 69 -3
rect 75 -9 81 -3
rect 87 -9 93 -3
rect 99 -9 105 -3
rect 111 -9 117 -3
rect 123 -9 129 -3
rect 135 -9 141 -3
rect 147 -9 153 -3
rect 159 -9 165 -3
rect 171 -9 177 -3
rect 183 -9 189 -3
rect 195 -9 201 -3
rect 207 -9 213 -3
rect 219 -9 225 -3
rect 231 -9 237 -3
rect 243 -9 249 -3
rect 255 -9 261 -3
rect 267 -9 273 -3
rect 279 -9 285 -3
rect 291 -9 297 -3
rect 303 -9 309 -3
rect 315 -9 321 -3
rect 327 -9 333 -3
rect 339 -9 345 -3
rect 351 -9 357 -3
rect 363 -9 369 -3
rect 375 -9 381 -3
rect 387 -9 393 -3
rect 399 -9 405 -3
rect 411 -9 417 -3
rect 423 -9 429 -3
rect 435 -9 441 -3
rect 447 -9 453 -3
rect 459 -9 465 -3
rect 471 -9 477 -3
rect 483 -9 489 -3
rect 495 -9 501 -3
rect 507 -9 513 -3
rect 519 -9 525 -3
rect 531 -9 537 -3
rect 543 -9 549 -3
rect 555 -9 561 -3
rect 567 -9 573 -3
rect 579 -9 585 -3
rect 591 -9 597 -3
rect 603 -9 609 -3
rect 615 -9 621 -3
rect 627 -9 633 -3
rect 639 -9 645 -3
rect 651 -9 657 -3
rect 663 -9 669 -3
rect 675 -9 681 -3
rect 687 -9 693 -3
rect 699 -9 705 -3
rect 711 -9 717 -3
rect 723 -9 729 -3
rect 735 -9 741 -3
rect 747 -9 753 -3
rect 759 -9 765 -3
rect 771 -9 777 -3
rect 783 -9 789 -3
rect 795 -9 801 -3
rect 807 -9 813 -3
rect 819 -9 825 -3
rect 831 -9 837 -3
rect 843 -9 849 -3
rect 855 -9 861 -3
rect 867 -9 873 -3
rect 879 -9 885 -3
rect 891 -9 897 -3
rect 903 -9 909 -3
rect 915 -9 921 -3
rect 927 -9 933 -3
rect 939 -9 945 -3
rect 951 -9 957 -3
rect 963 -9 969 -3
rect 975 -9 981 -3
rect 987 -9 993 -3
rect 999 -9 1005 -3
rect 1011 -9 1017 -3
rect 1023 -9 1029 -3
rect 1035 -9 1041 -3
rect 1047 -9 1053 -3
rect 1059 -9 1065 -3
rect 1071 -9 1077 -3
rect 1083 -9 1089 -3
rect 1095 -9 1101 -3
rect 1107 -9 1113 -3
rect 1119 -9 1125 -3
rect 1131 -9 1137 -3
rect 1143 -9 1149 -3
rect 1155 -9 1161 -3
rect 1167 -9 1173 -3
rect 1179 -9 1185 -3
rect 1191 -9 1197 -3
rect 1203 -9 1209 -3
rect 1215 -9 1221 -3
rect 1227 -9 1233 -3
rect 1239 -9 1245 -3
rect 1251 -9 1257 -3
rect 1263 -9 1269 -3
<< mvpsubdiffcont >>
rect -21 255 -15 261
rect -9 255 -3 261
rect 3 255 9 261
rect 15 255 21 261
rect 27 255 33 261
rect 39 255 45 261
rect 51 255 57 261
rect 63 255 69 261
rect 75 255 81 261
rect 87 255 93 261
rect 99 255 105 261
rect 111 255 117 261
rect 123 255 129 261
rect 135 255 141 261
rect 147 255 153 261
rect 159 255 165 261
rect 171 255 177 261
rect 183 255 189 261
rect 195 255 201 261
rect 207 255 213 261
rect 219 255 225 261
rect 231 255 237 261
rect 243 255 249 261
rect 255 255 261 261
rect 267 255 273 261
rect 279 255 285 261
rect 291 255 297 261
rect 303 255 309 261
rect 315 255 321 261
rect 327 255 333 261
rect 339 255 345 261
rect 351 255 357 261
rect 363 255 369 261
rect 375 255 381 261
rect 387 255 393 261
rect 399 255 405 261
rect 411 255 417 261
rect 423 255 429 261
rect 435 255 441 261
rect 447 255 453 261
rect 459 255 465 261
rect 471 255 477 261
rect 483 255 489 261
rect 495 255 501 261
rect 507 255 513 261
rect 519 255 525 261
rect 531 255 537 261
rect 543 255 549 261
rect 555 255 561 261
rect 567 255 573 261
rect 579 255 585 261
rect 591 255 597 261
rect 603 255 609 261
rect 615 255 621 261
rect 627 255 633 261
rect 639 255 645 261
rect 651 255 657 261
rect 663 255 669 261
rect 675 255 681 261
rect 687 255 693 261
rect 699 255 705 261
rect 711 255 717 261
rect 723 255 729 261
rect 735 255 741 261
rect 747 255 753 261
rect 759 255 765 261
rect 771 255 777 261
rect 783 255 789 261
rect 795 255 801 261
rect 807 255 813 261
rect 819 255 825 261
rect 831 255 837 261
rect 843 255 849 261
rect 855 255 861 261
rect 867 255 873 261
rect 879 255 885 261
rect 891 255 897 261
rect 903 255 909 261
rect 915 255 921 261
rect 927 255 933 261
rect 939 255 945 261
rect 951 255 957 261
rect 963 255 969 261
rect 975 255 981 261
rect 987 255 993 261
rect 999 255 1005 261
rect 1011 255 1017 261
rect 1023 255 1029 261
rect 1035 255 1041 261
rect 1047 255 1053 261
<< mvnsubdiffcont >>
rect -9 459 -3 465
rect 3 459 9 465
rect 15 459 21 465
rect 27 459 33 465
rect 39 459 45 465
rect 51 459 57 465
rect 63 459 69 465
rect 75 459 81 465
rect 87 459 93 465
rect 99 459 105 465
rect 111 459 117 465
rect 123 459 129 465
rect 135 459 141 465
rect 147 459 153 465
rect 159 459 165 465
rect 171 459 177 465
rect 183 459 189 465
rect 195 459 201 465
rect 207 459 213 465
rect 219 459 225 465
rect 231 459 237 465
rect 243 459 249 465
rect 255 459 261 465
rect 267 459 273 465
rect 279 459 285 465
rect 291 459 297 465
rect 303 459 309 465
rect 315 459 321 465
rect 327 459 333 465
rect 339 459 345 465
rect 351 459 357 465
rect 363 459 369 465
rect 375 459 381 465
rect 387 459 393 465
rect 399 459 405 465
rect 411 459 417 465
rect 423 459 429 465
rect 435 459 441 465
rect 447 459 453 465
rect 459 459 465 465
rect 471 459 477 465
rect 483 459 489 465
rect 495 459 501 465
rect 507 459 513 465
rect 519 459 525 465
rect 531 459 537 465
rect 543 459 549 465
rect 555 459 561 465
rect 567 459 573 465
rect 579 459 585 465
rect 591 459 597 465
rect 603 459 609 465
rect 615 459 621 465
rect 627 459 633 465
rect 639 459 645 465
rect 651 459 657 465
rect 663 459 669 465
rect 675 459 681 465
rect 687 459 693 465
rect 699 459 705 465
rect 711 459 717 465
rect 723 459 729 465
rect 735 459 741 465
rect 747 459 753 465
rect 759 459 765 465
rect 771 459 777 465
rect 783 459 789 465
rect 795 459 801 465
rect 807 459 813 465
rect 819 459 825 465
rect 831 459 837 465
rect 843 459 849 465
rect 855 459 861 465
rect 867 459 873 465
rect 879 459 885 465
rect 891 459 897 465
rect 903 459 909 465
rect 915 459 921 465
rect 927 459 933 465
rect 939 459 945 465
rect 951 459 957 465
rect 963 459 969 465
rect 975 459 981 465
rect 987 459 993 465
rect 999 459 1005 465
rect 1011 459 1017 465
rect 1023 459 1029 465
rect 1035 459 1041 465
rect 1047 459 1053 465
rect -9 279 -3 285
rect 3 279 9 285
rect 15 279 21 285
rect 27 279 33 285
rect 39 279 45 285
rect 51 279 57 285
rect 63 279 69 285
rect 75 279 81 285
rect 87 279 93 285
rect 99 279 105 285
rect 111 279 117 285
rect 123 279 129 285
rect 135 279 141 285
rect 147 279 153 285
rect 159 279 165 285
rect 171 279 177 285
rect 183 279 189 285
rect 195 279 201 285
rect 207 279 213 285
rect 219 279 225 285
rect 231 279 237 285
rect 243 279 249 285
rect 255 279 261 285
rect 267 279 273 285
rect 279 279 285 285
rect 291 279 297 285
rect 303 279 309 285
rect 315 279 321 285
rect 327 279 333 285
rect 339 279 345 285
rect 351 279 357 285
rect 363 279 369 285
rect 375 279 381 285
rect 387 279 393 285
rect 399 279 405 285
rect 411 279 417 285
rect 423 279 429 285
rect 435 279 441 285
rect 447 279 453 285
rect 459 279 465 285
rect 471 279 477 285
rect 483 279 489 285
rect 495 279 501 285
rect 507 279 513 285
rect 519 279 525 285
rect 531 279 537 285
rect 543 279 549 285
rect 555 279 561 285
rect 567 279 573 285
rect 579 279 585 285
rect 591 279 597 285
rect 603 279 609 285
rect 615 279 621 285
rect 627 279 633 285
rect 639 279 645 285
rect 651 279 657 285
rect 663 279 669 285
rect 675 279 681 285
rect 687 279 693 285
rect 699 279 705 285
rect 711 279 717 285
rect 723 279 729 285
rect 735 279 741 285
rect 747 279 753 285
rect 759 279 765 285
rect 771 279 777 285
rect 783 279 789 285
rect 795 279 801 285
rect 807 279 813 285
rect 819 279 825 285
rect 831 279 837 285
rect 843 279 849 285
rect 855 279 861 285
rect 867 279 873 285
rect 879 279 885 285
rect 891 279 897 285
rect 903 279 909 285
rect 915 279 921 285
rect 927 279 933 285
rect 939 279 945 285
rect 951 279 957 285
rect 963 279 969 285
rect 975 279 981 285
rect 987 279 993 285
rect 999 279 1005 285
rect 1011 279 1017 285
rect 1023 279 1029 285
rect 1035 279 1041 285
rect 1047 279 1053 285
<< polysilicon >>
rect 0 444 12 450
rect 24 444 36 450
rect 48 444 60 450
rect 72 444 84 450
rect 96 444 108 450
rect 120 444 132 450
rect 144 444 156 450
rect 168 444 180 450
rect 216 444 228 450
rect 240 444 252 450
rect 264 444 276 450
rect 288 444 300 450
rect 312 444 324 450
rect 336 444 348 450
rect 360 444 372 450
rect 384 444 396 450
rect 432 444 444 450
rect 456 444 468 450
rect 480 444 492 450
rect 504 444 516 450
rect 528 444 540 450
rect 552 444 564 450
rect 576 444 588 450
rect 600 444 612 450
rect 648 444 660 450
rect 672 444 684 450
rect 696 444 708 450
rect 720 444 732 450
rect 744 444 756 450
rect 768 444 780 450
rect 792 444 804 450
rect 816 444 828 450
rect 864 444 876 450
rect 888 444 900 450
rect 912 444 924 450
rect 936 444 948 450
rect 960 444 972 450
rect 984 444 996 450
rect 1008 444 1020 450
rect 1032 444 1044 450
rect 0 396 12 408
rect 24 396 36 408
rect 0 393 36 396
rect 0 387 3 393
rect 9 387 15 393
rect 21 387 27 393
rect 33 387 36 393
rect 0 384 36 387
rect 48 396 60 408
rect 72 396 84 408
rect 48 393 84 396
rect 48 387 51 393
rect 57 387 63 393
rect 69 387 75 393
rect 81 387 84 393
rect 48 384 84 387
rect 96 396 108 408
rect 120 396 132 408
rect 96 393 132 396
rect 96 387 99 393
rect 105 387 111 393
rect 117 387 123 393
rect 129 387 132 393
rect 96 384 132 387
rect 144 396 156 408
rect 168 396 180 408
rect 144 393 180 396
rect 144 387 147 393
rect 153 387 159 393
rect 165 387 171 393
rect 177 387 180 393
rect 144 384 180 387
rect 216 396 228 408
rect 240 396 252 408
rect 216 393 252 396
rect 216 387 219 393
rect 225 387 231 393
rect 237 387 243 393
rect 249 387 252 393
rect 216 384 252 387
rect 264 396 276 408
rect 288 396 300 408
rect 264 393 300 396
rect 264 387 267 393
rect 273 387 279 393
rect 285 387 291 393
rect 297 387 300 393
rect 264 384 300 387
rect 312 396 324 408
rect 336 396 348 408
rect 312 393 348 396
rect 312 387 315 393
rect 321 387 327 393
rect 333 387 339 393
rect 345 387 348 393
rect 312 384 348 387
rect 360 396 372 408
rect 384 396 396 408
rect 360 393 396 396
rect 360 387 363 393
rect 369 387 375 393
rect 381 387 387 393
rect 393 387 396 393
rect 360 384 396 387
rect 432 396 444 408
rect 456 396 468 408
rect 432 393 468 396
rect 432 387 435 393
rect 441 387 447 393
rect 453 387 459 393
rect 465 387 468 393
rect 432 384 468 387
rect 480 396 492 408
rect 504 396 516 408
rect 480 393 516 396
rect 480 387 483 393
rect 489 387 495 393
rect 501 387 507 393
rect 513 387 516 393
rect 480 384 516 387
rect 528 396 540 408
rect 552 396 564 408
rect 528 393 564 396
rect 528 387 531 393
rect 537 387 543 393
rect 549 387 555 393
rect 561 387 564 393
rect 528 384 564 387
rect 576 396 588 408
rect 600 396 612 408
rect 576 393 612 396
rect 576 387 579 393
rect 585 387 591 393
rect 597 387 603 393
rect 609 387 612 393
rect 576 384 612 387
rect 648 396 660 408
rect 672 396 684 408
rect 648 393 684 396
rect 648 387 651 393
rect 657 387 663 393
rect 669 387 675 393
rect 681 387 684 393
rect 648 384 684 387
rect 696 396 708 408
rect 720 396 732 408
rect 696 393 732 396
rect 696 387 699 393
rect 705 387 711 393
rect 717 387 723 393
rect 729 387 732 393
rect 696 384 732 387
rect 744 396 756 408
rect 768 396 780 408
rect 744 393 780 396
rect 744 387 747 393
rect 753 387 759 393
rect 765 387 771 393
rect 777 387 780 393
rect 744 384 780 387
rect 792 396 804 408
rect 816 396 828 408
rect 792 393 828 396
rect 792 387 795 393
rect 801 387 807 393
rect 813 387 819 393
rect 825 387 828 393
rect 792 384 828 387
rect 864 396 876 408
rect 888 396 900 408
rect 912 396 924 408
rect 936 396 948 408
rect 864 393 948 396
rect 864 387 867 393
rect 873 387 879 393
rect 885 387 891 393
rect 897 387 903 393
rect 909 387 915 393
rect 921 387 927 393
rect 933 387 939 393
rect 945 387 948 393
rect 864 384 948 387
rect 960 396 972 408
rect 984 396 996 408
rect 960 393 996 396
rect 960 387 963 393
rect 969 387 975 393
rect 981 387 987 393
rect 993 387 996 393
rect 960 384 996 387
rect 1008 396 1020 408
rect 1032 396 1044 408
rect 1008 393 1044 396
rect 1008 387 1011 393
rect 1017 387 1023 393
rect 1029 387 1035 393
rect 1041 387 1044 393
rect 1008 384 1044 387
rect 0 360 12 366
rect 24 360 36 366
rect 48 360 60 366
rect 72 360 84 366
rect 96 360 108 366
rect 120 360 132 366
rect 144 360 156 366
rect 168 360 180 366
rect 216 360 228 366
rect 240 360 252 366
rect 264 360 276 366
rect 288 360 300 366
rect 312 360 324 366
rect 336 360 348 366
rect 360 360 372 366
rect 384 360 396 366
rect 432 360 444 366
rect 456 360 468 366
rect 480 360 492 366
rect 504 360 516 366
rect 528 360 540 366
rect 552 360 564 366
rect 576 360 588 366
rect 600 360 612 366
rect 648 360 660 366
rect 672 360 684 366
rect 696 360 708 366
rect 720 360 732 366
rect 744 360 756 366
rect 768 360 780 366
rect 792 360 804 366
rect 816 360 828 366
rect 864 360 876 366
rect 888 360 900 366
rect 912 360 924 366
rect 936 360 948 366
rect 960 360 972 366
rect 984 360 996 366
rect 1008 360 1020 366
rect 1032 360 1044 366
rect 0 312 12 324
rect 24 312 36 324
rect 0 309 36 312
rect 0 303 3 309
rect 9 303 15 309
rect 21 303 27 309
rect 33 303 36 309
rect 0 300 36 303
rect 48 312 60 324
rect 72 312 84 324
rect 48 309 84 312
rect 48 303 51 309
rect 57 303 63 309
rect 69 303 75 309
rect 81 303 84 309
rect 48 300 84 303
rect 96 312 108 324
rect 120 312 132 324
rect 96 309 132 312
rect 96 303 99 309
rect 105 303 111 309
rect 117 303 123 309
rect 129 303 132 309
rect 96 300 132 303
rect 144 312 156 324
rect 168 312 180 324
rect 144 309 180 312
rect 144 303 147 309
rect 153 303 159 309
rect 165 303 171 309
rect 177 303 180 309
rect 144 300 180 303
rect 216 312 228 324
rect 240 312 252 324
rect 216 309 252 312
rect 216 303 219 309
rect 225 303 231 309
rect 237 303 243 309
rect 249 303 252 309
rect 216 300 252 303
rect 264 312 276 324
rect 288 312 300 324
rect 264 309 300 312
rect 264 303 267 309
rect 273 303 279 309
rect 285 303 291 309
rect 297 303 300 309
rect 264 300 300 303
rect 312 312 324 324
rect 336 312 348 324
rect 312 309 348 312
rect 312 303 315 309
rect 321 303 327 309
rect 333 303 339 309
rect 345 303 348 309
rect 312 300 348 303
rect 360 312 372 324
rect 384 312 396 324
rect 360 309 396 312
rect 360 303 363 309
rect 369 303 375 309
rect 381 303 387 309
rect 393 303 396 309
rect 360 300 396 303
rect 432 312 444 324
rect 456 312 468 324
rect 432 309 468 312
rect 432 303 435 309
rect 441 303 447 309
rect 453 303 459 309
rect 465 303 468 309
rect 432 300 468 303
rect 480 312 492 324
rect 504 312 516 324
rect 480 309 516 312
rect 480 303 483 309
rect 489 303 495 309
rect 501 303 507 309
rect 513 303 516 309
rect 480 300 516 303
rect 528 312 540 324
rect 552 312 564 324
rect 528 309 564 312
rect 528 303 531 309
rect 537 303 543 309
rect 549 303 555 309
rect 561 303 564 309
rect 528 300 564 303
rect 576 312 588 324
rect 600 312 612 324
rect 576 309 612 312
rect 576 303 579 309
rect 585 303 591 309
rect 597 303 603 309
rect 609 303 612 309
rect 576 300 612 303
rect 648 312 660 324
rect 672 312 684 324
rect 648 309 684 312
rect 648 303 651 309
rect 657 303 663 309
rect 669 303 675 309
rect 681 303 684 309
rect 648 300 684 303
rect 696 312 708 324
rect 720 312 732 324
rect 696 309 732 312
rect 696 303 699 309
rect 705 303 711 309
rect 717 303 723 309
rect 729 303 732 309
rect 696 300 732 303
rect 744 312 756 324
rect 768 312 780 324
rect 744 309 780 312
rect 744 303 747 309
rect 753 303 759 309
rect 765 303 771 309
rect 777 303 780 309
rect 744 300 780 303
rect 792 312 804 324
rect 816 312 828 324
rect 792 309 828 312
rect 792 303 795 309
rect 801 303 807 309
rect 813 303 819 309
rect 825 303 828 309
rect 792 300 828 303
rect 864 312 876 324
rect 888 312 900 324
rect 912 312 924 324
rect 936 312 948 324
rect 864 309 948 312
rect 864 303 867 309
rect 873 303 879 309
rect 885 303 891 309
rect 897 303 903 309
rect 909 303 915 309
rect 921 303 927 309
rect 933 303 939 309
rect 945 303 948 309
rect 864 300 948 303
rect 960 312 972 324
rect 984 312 996 324
rect 960 309 996 312
rect 960 303 963 309
rect 969 303 975 309
rect 981 303 987 309
rect 993 303 996 309
rect 960 300 996 303
rect 1008 312 1020 324
rect 1032 312 1044 324
rect 1008 309 1044 312
rect 1008 303 1011 309
rect 1017 303 1023 309
rect 1029 303 1035 309
rect 1041 303 1044 309
rect 1008 300 1044 303
rect 0 237 36 240
rect 0 231 3 237
rect 9 231 15 237
rect 21 231 27 237
rect 33 231 36 237
rect 0 228 36 231
rect 0 216 12 228
rect 24 216 36 228
rect 48 237 84 240
rect 48 231 51 237
rect 57 231 63 237
rect 69 231 75 237
rect 81 231 84 237
rect 48 228 84 231
rect 48 216 60 228
rect 72 216 84 228
rect 96 237 132 240
rect 96 231 99 237
rect 105 231 111 237
rect 117 231 123 237
rect 129 231 132 237
rect 96 228 132 231
rect 96 216 108 228
rect 120 216 132 228
rect 144 237 180 240
rect 144 231 147 237
rect 153 231 159 237
rect 165 231 171 237
rect 177 231 180 237
rect 144 228 180 231
rect 144 216 156 228
rect 168 216 180 228
rect 216 237 252 240
rect 216 231 219 237
rect 225 231 231 237
rect 237 231 243 237
rect 249 231 252 237
rect 216 228 252 231
rect 216 216 228 228
rect 240 216 252 228
rect 264 237 300 240
rect 264 231 267 237
rect 273 231 279 237
rect 285 231 291 237
rect 297 231 300 237
rect 264 228 300 231
rect 264 216 276 228
rect 288 216 300 228
rect 312 237 348 240
rect 312 231 315 237
rect 321 231 327 237
rect 333 231 339 237
rect 345 231 348 237
rect 312 228 348 231
rect 312 216 324 228
rect 336 216 348 228
rect 360 237 396 240
rect 360 231 363 237
rect 369 231 375 237
rect 381 231 387 237
rect 393 231 396 237
rect 360 228 396 231
rect 360 216 372 228
rect 384 216 396 228
rect 432 237 468 240
rect 432 231 435 237
rect 441 231 447 237
rect 453 231 459 237
rect 465 231 468 237
rect 432 228 468 231
rect 432 216 444 228
rect 456 216 468 228
rect 480 237 516 240
rect 480 231 483 237
rect 489 231 495 237
rect 501 231 507 237
rect 513 231 516 237
rect 480 228 516 231
rect 480 216 492 228
rect 504 216 516 228
rect 528 237 564 240
rect 528 231 531 237
rect 537 231 543 237
rect 549 231 555 237
rect 561 231 564 237
rect 528 228 564 231
rect 528 216 540 228
rect 552 216 564 228
rect 576 237 612 240
rect 576 231 579 237
rect 585 231 591 237
rect 597 231 603 237
rect 609 231 612 237
rect 576 228 612 231
rect 576 216 588 228
rect 600 216 612 228
rect 648 237 684 240
rect 648 231 651 237
rect 657 231 663 237
rect 669 231 675 237
rect 681 231 684 237
rect 648 228 684 231
rect 648 216 660 228
rect 672 216 684 228
rect 696 237 732 240
rect 696 231 699 237
rect 705 231 711 237
rect 717 231 723 237
rect 729 231 732 237
rect 696 228 732 231
rect 696 216 708 228
rect 720 216 732 228
rect 744 237 780 240
rect 744 231 747 237
rect 753 231 759 237
rect 765 231 771 237
rect 777 231 780 237
rect 744 228 780 231
rect 744 216 756 228
rect 768 216 780 228
rect 792 237 828 240
rect 792 231 795 237
rect 801 231 807 237
rect 813 231 819 237
rect 825 231 828 237
rect 792 228 828 231
rect 792 216 804 228
rect 816 216 828 228
rect 864 237 876 240
rect 864 231 867 237
rect 873 231 876 237
rect 864 216 876 231
rect 912 237 948 240
rect 912 231 915 237
rect 921 231 927 237
rect 933 231 939 237
rect 945 231 948 237
rect 912 228 948 231
rect 912 216 924 228
rect 936 216 948 228
rect 960 237 996 240
rect 960 231 963 237
rect 969 231 975 237
rect 981 231 987 237
rect 993 231 996 237
rect 960 228 996 231
rect 960 216 972 228
rect 984 216 996 228
rect 1008 237 1044 240
rect 1008 231 1011 237
rect 1017 231 1023 237
rect 1029 231 1035 237
rect 1041 231 1044 237
rect 1008 228 1044 231
rect 1008 216 1020 228
rect 1032 216 1044 228
rect 1080 237 1116 240
rect 1080 231 1083 237
rect 1089 231 1095 237
rect 1101 231 1107 237
rect 1113 231 1116 237
rect 1080 228 1116 231
rect 1080 216 1092 228
rect 1104 216 1116 228
rect 1128 237 1164 240
rect 1128 231 1131 237
rect 1137 231 1143 237
rect 1149 231 1155 237
rect 1161 231 1164 237
rect 1128 228 1164 231
rect 1128 216 1140 228
rect 1152 216 1164 228
rect 1176 237 1212 240
rect 1176 231 1179 237
rect 1185 231 1191 237
rect 1197 231 1203 237
rect 1209 231 1212 237
rect 1176 228 1212 231
rect 1176 216 1188 228
rect 1200 216 1212 228
rect 1224 237 1260 240
rect 1224 231 1227 237
rect 1233 231 1239 237
rect 1245 231 1251 237
rect 1257 231 1260 237
rect 1224 228 1260 231
rect 1224 216 1236 228
rect 1248 216 1260 228
rect 0 174 12 180
rect 24 174 36 180
rect 48 174 60 180
rect 72 174 84 180
rect 96 174 108 180
rect 120 174 132 180
rect 144 174 156 180
rect 168 174 180 180
rect 216 174 228 180
rect 240 174 252 180
rect 264 174 276 180
rect 288 174 300 180
rect 312 174 324 180
rect 336 174 348 180
rect 360 174 372 180
rect 384 174 396 180
rect 432 174 444 180
rect 456 174 468 180
rect 480 174 492 180
rect 504 174 516 180
rect 528 174 540 180
rect 552 174 564 180
rect 576 174 588 180
rect 600 174 612 180
rect 648 174 660 180
rect 672 174 684 180
rect 696 174 708 180
rect 720 174 732 180
rect 744 174 756 180
rect 768 174 780 180
rect 792 174 804 180
rect 816 174 828 180
rect 864 174 876 180
rect 912 174 924 180
rect 936 174 948 180
rect 960 174 972 180
rect 984 174 996 180
rect 1008 174 1020 180
rect 1032 174 1044 180
rect 1080 174 1092 180
rect 1104 174 1116 180
rect 1128 174 1140 180
rect 1152 174 1164 180
rect 1176 174 1188 180
rect 1200 174 1212 180
rect 1224 174 1236 180
rect 1248 174 1260 180
rect 0 69 36 72
rect 0 63 3 69
rect 9 63 15 69
rect 21 63 27 69
rect 33 63 36 69
rect 0 60 36 63
rect 0 48 12 60
rect 24 48 36 60
rect 48 69 84 72
rect 48 63 51 69
rect 57 63 63 69
rect 69 63 75 69
rect 81 63 84 69
rect 48 60 84 63
rect 48 48 60 60
rect 72 48 84 60
rect 96 69 132 72
rect 96 63 99 69
rect 105 63 111 69
rect 117 63 123 69
rect 129 63 132 69
rect 96 60 132 63
rect 96 48 108 60
rect 120 48 132 60
rect 144 69 180 72
rect 144 63 147 69
rect 153 63 159 69
rect 165 63 171 69
rect 177 63 180 69
rect 144 60 180 63
rect 144 48 156 60
rect 168 48 180 60
rect 216 69 252 72
rect 216 63 219 69
rect 225 63 231 69
rect 237 63 243 69
rect 249 63 252 69
rect 216 60 252 63
rect 216 48 228 60
rect 240 48 252 60
rect 264 69 300 72
rect 264 63 267 69
rect 273 63 279 69
rect 285 63 291 69
rect 297 63 300 69
rect 264 60 300 63
rect 264 48 276 60
rect 288 48 300 60
rect 312 69 348 72
rect 312 63 315 69
rect 321 63 327 69
rect 333 63 339 69
rect 345 63 348 69
rect 312 60 348 63
rect 312 48 324 60
rect 336 48 348 60
rect 360 69 396 72
rect 360 63 363 69
rect 369 63 375 69
rect 381 63 387 69
rect 393 63 396 69
rect 360 60 396 63
rect 360 48 372 60
rect 384 48 396 60
rect 432 69 468 72
rect 432 63 435 69
rect 441 63 447 69
rect 453 63 459 69
rect 465 63 468 69
rect 432 60 468 63
rect 432 48 444 60
rect 456 48 468 60
rect 480 69 516 72
rect 480 63 483 69
rect 489 63 495 69
rect 501 63 507 69
rect 513 63 516 69
rect 480 60 516 63
rect 480 48 492 60
rect 504 48 516 60
rect 528 69 564 72
rect 528 63 531 69
rect 537 63 543 69
rect 549 63 555 69
rect 561 63 564 69
rect 528 60 564 63
rect 528 48 540 60
rect 552 48 564 60
rect 576 69 612 72
rect 576 63 579 69
rect 585 63 591 69
rect 597 63 603 69
rect 609 63 612 69
rect 576 60 612 63
rect 576 48 588 60
rect 600 48 612 60
rect 648 69 684 72
rect 648 63 651 69
rect 657 63 663 69
rect 669 63 675 69
rect 681 63 684 69
rect 648 60 684 63
rect 648 48 660 60
rect 672 48 684 60
rect 696 69 732 72
rect 696 63 699 69
rect 705 63 711 69
rect 717 63 723 69
rect 729 63 732 69
rect 696 60 732 63
rect 696 48 708 60
rect 720 48 732 60
rect 744 69 780 72
rect 744 63 747 69
rect 753 63 759 69
rect 765 63 771 69
rect 777 63 780 69
rect 744 60 780 63
rect 744 48 756 60
rect 768 48 780 60
rect 792 69 828 72
rect 792 63 795 69
rect 801 63 807 69
rect 813 63 819 69
rect 825 63 828 69
rect 792 60 828 63
rect 792 48 804 60
rect 816 48 828 60
rect 864 69 900 72
rect 864 63 867 69
rect 873 63 879 69
rect 885 63 891 69
rect 897 63 900 69
rect 864 60 900 63
rect 864 48 876 60
rect 888 48 900 60
rect 912 69 948 72
rect 912 63 915 69
rect 921 63 927 69
rect 933 63 939 69
rect 945 63 948 69
rect 912 60 948 63
rect 912 48 924 60
rect 936 48 948 60
rect 960 69 996 72
rect 960 63 963 69
rect 969 63 975 69
rect 981 63 987 69
rect 993 63 996 69
rect 960 60 996 63
rect 960 48 972 60
rect 984 48 996 60
rect 1008 69 1044 72
rect 1008 63 1011 69
rect 1017 63 1023 69
rect 1029 63 1035 69
rect 1041 63 1044 69
rect 1008 60 1044 63
rect 1008 48 1020 60
rect 1032 48 1044 60
rect 1080 69 1116 72
rect 1080 63 1083 69
rect 1089 63 1095 69
rect 1101 63 1107 69
rect 1113 63 1116 69
rect 1080 60 1116 63
rect 1080 48 1092 60
rect 1104 48 1116 60
rect 1128 69 1164 72
rect 1128 63 1131 69
rect 1137 63 1143 69
rect 1149 63 1155 69
rect 1161 63 1164 69
rect 1128 60 1164 63
rect 1128 48 1140 60
rect 1152 48 1164 60
rect 1176 69 1212 72
rect 1176 63 1179 69
rect 1185 63 1191 69
rect 1197 63 1203 69
rect 1209 63 1212 69
rect 1176 60 1212 63
rect 1176 48 1188 60
rect 1200 48 1212 60
rect 1224 69 1260 72
rect 1224 63 1227 69
rect 1233 63 1239 69
rect 1245 63 1251 69
rect 1257 63 1260 69
rect 1224 60 1260 63
rect 1224 48 1236 60
rect 1248 48 1260 60
rect 0 6 12 12
rect 24 6 36 12
rect 48 6 60 12
rect 72 6 84 12
rect 96 6 108 12
rect 120 6 132 12
rect 144 6 156 12
rect 168 6 180 12
rect 216 6 228 12
rect 240 6 252 12
rect 264 6 276 12
rect 288 6 300 12
rect 312 6 324 12
rect 336 6 348 12
rect 360 6 372 12
rect 384 6 396 12
rect 432 6 444 12
rect 456 6 468 12
rect 480 6 492 12
rect 504 6 516 12
rect 528 6 540 12
rect 552 6 564 12
rect 576 6 588 12
rect 600 6 612 12
rect 648 6 660 12
rect 672 6 684 12
rect 696 6 708 12
rect 720 6 732 12
rect 744 6 756 12
rect 768 6 780 12
rect 792 6 804 12
rect 816 6 828 12
rect 864 6 876 12
rect 888 6 900 12
rect 912 6 924 12
rect 936 6 948 12
rect 960 6 972 12
rect 984 6 996 12
rect 1008 6 1020 12
rect 1032 6 1044 12
rect 1080 6 1092 12
rect 1104 6 1116 12
rect 1128 6 1140 12
rect 1152 6 1164 12
rect 1176 6 1188 12
rect 1200 6 1212 12
rect 1224 6 1236 12
rect 1248 6 1260 12
<< polycontact >>
rect 3 387 9 393
rect 15 387 21 393
rect 27 387 33 393
rect 51 387 57 393
rect 63 387 69 393
rect 75 387 81 393
rect 99 387 105 393
rect 111 387 117 393
rect 123 387 129 393
rect 147 387 153 393
rect 159 387 165 393
rect 171 387 177 393
rect 219 387 225 393
rect 231 387 237 393
rect 243 387 249 393
rect 267 387 273 393
rect 279 387 285 393
rect 291 387 297 393
rect 315 387 321 393
rect 327 387 333 393
rect 339 387 345 393
rect 363 387 369 393
rect 375 387 381 393
rect 387 387 393 393
rect 435 387 441 393
rect 447 387 453 393
rect 459 387 465 393
rect 483 387 489 393
rect 495 387 501 393
rect 507 387 513 393
rect 531 387 537 393
rect 543 387 549 393
rect 555 387 561 393
rect 579 387 585 393
rect 591 387 597 393
rect 603 387 609 393
rect 651 387 657 393
rect 663 387 669 393
rect 675 387 681 393
rect 699 387 705 393
rect 711 387 717 393
rect 723 387 729 393
rect 747 387 753 393
rect 759 387 765 393
rect 771 387 777 393
rect 795 387 801 393
rect 807 387 813 393
rect 819 387 825 393
rect 867 387 873 393
rect 879 387 885 393
rect 891 387 897 393
rect 903 387 909 393
rect 915 387 921 393
rect 927 387 933 393
rect 939 387 945 393
rect 963 387 969 393
rect 975 387 981 393
rect 987 387 993 393
rect 1011 387 1017 393
rect 1023 387 1029 393
rect 1035 387 1041 393
rect 3 303 9 309
rect 15 303 21 309
rect 27 303 33 309
rect 51 303 57 309
rect 63 303 69 309
rect 75 303 81 309
rect 99 303 105 309
rect 111 303 117 309
rect 123 303 129 309
rect 147 303 153 309
rect 159 303 165 309
rect 171 303 177 309
rect 219 303 225 309
rect 231 303 237 309
rect 243 303 249 309
rect 267 303 273 309
rect 279 303 285 309
rect 291 303 297 309
rect 315 303 321 309
rect 327 303 333 309
rect 339 303 345 309
rect 363 303 369 309
rect 375 303 381 309
rect 387 303 393 309
rect 435 303 441 309
rect 447 303 453 309
rect 459 303 465 309
rect 483 303 489 309
rect 495 303 501 309
rect 507 303 513 309
rect 531 303 537 309
rect 543 303 549 309
rect 555 303 561 309
rect 579 303 585 309
rect 591 303 597 309
rect 603 303 609 309
rect 651 303 657 309
rect 663 303 669 309
rect 675 303 681 309
rect 699 303 705 309
rect 711 303 717 309
rect 723 303 729 309
rect 747 303 753 309
rect 759 303 765 309
rect 771 303 777 309
rect 795 303 801 309
rect 807 303 813 309
rect 819 303 825 309
rect 867 303 873 309
rect 879 303 885 309
rect 891 303 897 309
rect 903 303 909 309
rect 915 303 921 309
rect 927 303 933 309
rect 939 303 945 309
rect 963 303 969 309
rect 975 303 981 309
rect 987 303 993 309
rect 1011 303 1017 309
rect 1023 303 1029 309
rect 1035 303 1041 309
rect 3 231 9 237
rect 15 231 21 237
rect 27 231 33 237
rect 51 231 57 237
rect 63 231 69 237
rect 75 231 81 237
rect 99 231 105 237
rect 111 231 117 237
rect 123 231 129 237
rect 147 231 153 237
rect 159 231 165 237
rect 171 231 177 237
rect 219 231 225 237
rect 231 231 237 237
rect 243 231 249 237
rect 267 231 273 237
rect 279 231 285 237
rect 291 231 297 237
rect 315 231 321 237
rect 327 231 333 237
rect 339 231 345 237
rect 363 231 369 237
rect 375 231 381 237
rect 387 231 393 237
rect 435 231 441 237
rect 447 231 453 237
rect 459 231 465 237
rect 483 231 489 237
rect 495 231 501 237
rect 507 231 513 237
rect 531 231 537 237
rect 543 231 549 237
rect 555 231 561 237
rect 579 231 585 237
rect 591 231 597 237
rect 603 231 609 237
rect 651 231 657 237
rect 663 231 669 237
rect 675 231 681 237
rect 699 231 705 237
rect 711 231 717 237
rect 723 231 729 237
rect 747 231 753 237
rect 759 231 765 237
rect 771 231 777 237
rect 795 231 801 237
rect 807 231 813 237
rect 819 231 825 237
rect 867 231 873 237
rect 915 231 921 237
rect 927 231 933 237
rect 939 231 945 237
rect 963 231 969 237
rect 975 231 981 237
rect 987 231 993 237
rect 1011 231 1017 237
rect 1023 231 1029 237
rect 1035 231 1041 237
rect 1083 231 1089 237
rect 1095 231 1101 237
rect 1107 231 1113 237
rect 1131 231 1137 237
rect 1143 231 1149 237
rect 1155 231 1161 237
rect 1179 231 1185 237
rect 1191 231 1197 237
rect 1203 231 1209 237
rect 1227 231 1233 237
rect 1239 231 1245 237
rect 1251 231 1257 237
rect 3 63 9 69
rect 15 63 21 69
rect 27 63 33 69
rect 51 63 57 69
rect 63 63 69 69
rect 75 63 81 69
rect 99 63 105 69
rect 111 63 117 69
rect 123 63 129 69
rect 147 63 153 69
rect 159 63 165 69
rect 171 63 177 69
rect 219 63 225 69
rect 231 63 237 69
rect 243 63 249 69
rect 267 63 273 69
rect 279 63 285 69
rect 291 63 297 69
rect 315 63 321 69
rect 327 63 333 69
rect 339 63 345 69
rect 363 63 369 69
rect 375 63 381 69
rect 387 63 393 69
rect 435 63 441 69
rect 447 63 453 69
rect 459 63 465 69
rect 483 63 489 69
rect 495 63 501 69
rect 507 63 513 69
rect 531 63 537 69
rect 543 63 549 69
rect 555 63 561 69
rect 579 63 585 69
rect 591 63 597 69
rect 603 63 609 69
rect 651 63 657 69
rect 663 63 669 69
rect 675 63 681 69
rect 699 63 705 69
rect 711 63 717 69
rect 723 63 729 69
rect 747 63 753 69
rect 759 63 765 69
rect 771 63 777 69
rect 795 63 801 69
rect 807 63 813 69
rect 819 63 825 69
rect 867 63 873 69
rect 879 63 885 69
rect 891 63 897 69
rect 915 63 921 69
rect 927 63 933 69
rect 939 63 945 69
rect 963 63 969 69
rect 975 63 981 69
rect 987 63 993 69
rect 1011 63 1017 69
rect 1023 63 1029 69
rect 1035 63 1041 69
rect 1083 63 1089 69
rect 1095 63 1101 69
rect 1107 63 1113 69
rect 1131 63 1137 69
rect 1143 63 1149 69
rect 1155 63 1161 69
rect 1179 63 1185 69
rect 1191 63 1197 69
rect 1203 63 1209 69
rect 1227 63 1233 69
rect 1239 63 1245 69
rect 1251 63 1257 69
<< metal1 >>
rect -12 465 1056 468
rect -12 459 -9 465
rect -3 459 3 465
rect 9 459 15 465
rect 21 459 27 465
rect 33 459 39 465
rect 45 459 51 465
rect 57 459 63 465
rect 69 459 75 465
rect 81 459 87 465
rect 93 459 99 465
rect 105 459 111 465
rect 117 459 123 465
rect 129 459 135 465
rect 141 459 147 465
rect 153 459 159 465
rect 165 459 171 465
rect 177 459 183 465
rect 189 459 195 465
rect 201 459 207 465
rect 213 459 219 465
rect 225 459 231 465
rect 237 459 243 465
rect 249 459 255 465
rect 261 459 267 465
rect 273 459 279 465
rect 285 459 291 465
rect 297 459 303 465
rect 309 459 315 465
rect 321 459 327 465
rect 333 459 339 465
rect 345 459 351 465
rect 357 459 363 465
rect 369 459 375 465
rect 381 459 387 465
rect 393 459 399 465
rect 405 459 411 465
rect 417 459 423 465
rect 429 459 435 465
rect 441 459 447 465
rect 453 459 459 465
rect 465 459 471 465
rect 477 459 483 465
rect 489 459 495 465
rect 501 459 507 465
rect 513 459 519 465
rect 525 459 531 465
rect 537 459 543 465
rect 549 459 555 465
rect 561 459 567 465
rect 573 459 579 465
rect 585 459 591 465
rect 597 459 603 465
rect 609 459 615 465
rect 621 459 627 465
rect 633 459 639 465
rect 645 459 651 465
rect 657 459 663 465
rect 669 459 675 465
rect 681 459 687 465
rect 693 459 699 465
rect 705 459 711 465
rect 717 459 723 465
rect 729 459 735 465
rect 741 459 747 465
rect 753 459 759 465
rect 765 459 771 465
rect 777 459 783 465
rect 789 459 795 465
rect 801 459 807 465
rect 813 459 819 465
rect 825 459 831 465
rect 837 459 843 465
rect 849 459 855 465
rect 861 459 867 465
rect 873 459 879 465
rect 885 459 891 465
rect 897 459 903 465
rect 909 459 915 465
rect 921 459 927 465
rect 933 459 939 465
rect 945 459 951 465
rect 957 459 963 465
rect 969 459 975 465
rect 981 459 987 465
rect 993 459 999 465
rect 1005 459 1011 465
rect 1017 459 1023 465
rect 1029 459 1035 465
rect 1041 459 1047 465
rect 1053 459 1056 465
rect -12 456 1056 459
rect -12 441 0 456
rect -12 435 -9 441
rect -3 435 0 441
rect -12 429 0 435
rect -12 423 -9 429
rect -3 423 0 429
rect -12 417 0 423
rect -12 411 -9 417
rect -3 411 0 417
rect -12 408 0 411
rect 12 441 24 444
rect 12 435 15 441
rect 21 435 24 441
rect 12 429 24 435
rect 12 423 15 429
rect 21 423 24 429
rect 12 417 24 423
rect 12 411 15 417
rect 21 411 24 417
rect 12 408 24 411
rect 36 441 48 456
rect 36 435 39 441
rect 45 435 48 441
rect 36 429 48 435
rect 36 423 39 429
rect 45 423 48 429
rect 36 417 48 423
rect 36 411 39 417
rect 45 411 48 417
rect 36 408 48 411
rect 60 441 72 444
rect 60 435 63 441
rect 69 435 72 441
rect 60 429 72 435
rect 60 423 63 429
rect 69 423 72 429
rect 60 417 72 423
rect 60 411 63 417
rect 69 411 72 417
rect 60 408 72 411
rect 84 441 96 456
rect 84 435 87 441
rect 93 435 96 441
rect 84 429 96 435
rect 84 423 87 429
rect 93 423 96 429
rect 84 417 96 423
rect 84 411 87 417
rect 93 411 96 417
rect 84 408 96 411
rect 108 441 120 444
rect 108 435 111 441
rect 117 435 120 441
rect 108 429 120 435
rect 108 423 111 429
rect 117 423 120 429
rect 108 417 120 423
rect 108 411 111 417
rect 117 411 120 417
rect 108 408 120 411
rect 132 441 144 456
rect 132 435 135 441
rect 141 435 144 441
rect 132 429 144 435
rect 132 423 135 429
rect 141 423 144 429
rect 132 417 144 423
rect 132 411 135 417
rect 141 411 144 417
rect 132 408 144 411
rect 156 441 168 444
rect 156 435 159 441
rect 165 435 168 441
rect 156 429 168 435
rect 156 423 159 429
rect 165 423 168 429
rect 156 417 168 423
rect 156 411 159 417
rect 165 411 168 417
rect 156 408 168 411
rect 180 441 192 456
rect 180 435 183 441
rect 189 435 192 441
rect 180 429 192 435
rect 180 423 183 429
rect 189 423 192 429
rect 180 417 192 423
rect 180 411 183 417
rect 189 411 192 417
rect 180 408 192 411
rect 204 441 216 456
rect 204 435 207 441
rect 213 435 216 441
rect 204 429 216 435
rect 204 423 207 429
rect 213 423 216 429
rect 204 417 216 423
rect 204 411 207 417
rect 213 411 216 417
rect 204 408 216 411
rect 252 441 264 444
rect 252 435 255 441
rect 261 435 264 441
rect 252 429 264 435
rect 252 423 255 429
rect 261 423 264 429
rect 252 417 264 423
rect 252 411 255 417
rect 261 411 264 417
rect 252 408 264 411
rect 300 441 312 456
rect 300 435 303 441
rect 309 435 312 441
rect 300 429 312 435
rect 300 423 303 429
rect 309 423 312 429
rect 300 417 312 423
rect 300 411 303 417
rect 309 411 312 417
rect 300 408 312 411
rect 348 441 360 444
rect 348 435 351 441
rect 357 435 360 441
rect 348 429 360 435
rect 348 423 351 429
rect 357 423 360 429
rect 348 417 360 423
rect 348 411 351 417
rect 357 411 360 417
rect 348 408 360 411
rect 396 441 408 456
rect 396 435 399 441
rect 405 435 408 441
rect 396 429 408 435
rect 396 423 399 429
rect 405 423 408 429
rect 396 417 408 423
rect 396 411 399 417
rect 405 411 408 417
rect 396 408 408 411
rect 420 441 432 456
rect 420 435 423 441
rect 429 435 432 441
rect 420 429 432 435
rect 420 423 423 429
rect 429 423 432 429
rect 420 417 432 423
rect 420 411 423 417
rect 429 411 432 417
rect 420 408 432 411
rect 468 441 480 444
rect 468 435 471 441
rect 477 435 480 441
rect 468 429 480 435
rect 468 423 471 429
rect 477 423 480 429
rect 468 417 480 423
rect 468 411 471 417
rect 477 411 480 417
rect 468 408 480 411
rect 516 441 528 456
rect 516 435 519 441
rect 525 435 528 441
rect 516 429 528 435
rect 516 423 519 429
rect 525 423 528 429
rect 516 417 528 423
rect 516 411 519 417
rect 525 411 528 417
rect 516 408 528 411
rect 564 441 576 444
rect 564 435 567 441
rect 573 435 576 441
rect 564 429 576 435
rect 564 423 567 429
rect 573 423 576 429
rect 564 417 576 423
rect 564 411 567 417
rect 573 411 576 417
rect 564 408 576 411
rect 612 441 624 456
rect 612 435 615 441
rect 621 435 624 441
rect 612 429 624 435
rect 612 423 615 429
rect 621 423 624 429
rect 612 417 624 423
rect 612 411 615 417
rect 621 411 624 417
rect 612 408 624 411
rect 636 441 648 456
rect 636 435 639 441
rect 645 435 648 441
rect 636 429 648 435
rect 636 423 639 429
rect 645 423 648 429
rect 636 417 648 423
rect 636 411 639 417
rect 645 411 648 417
rect 636 408 648 411
rect 828 441 840 444
rect 828 435 831 441
rect 837 435 840 441
rect 828 429 840 435
rect 828 423 831 429
rect 837 423 840 429
rect 828 417 840 423
rect 828 411 831 417
rect 837 411 840 417
rect 828 408 840 411
rect 852 441 864 456
rect 852 435 855 441
rect 861 435 864 441
rect 852 429 864 435
rect 852 423 855 429
rect 861 423 864 429
rect 852 417 864 423
rect 852 411 855 417
rect 861 411 864 417
rect 852 408 864 411
rect 1044 441 1056 444
rect 1044 435 1047 441
rect 1053 435 1056 441
rect 1044 429 1056 435
rect 1044 423 1047 429
rect 1053 423 1056 429
rect 1044 417 1056 423
rect 1044 411 1047 417
rect 1053 411 1056 417
rect 1044 408 1056 411
rect 0 393 180 396
rect 0 387 3 393
rect 9 387 15 393
rect 21 387 27 393
rect 33 387 39 393
rect 45 387 51 393
rect 57 387 63 393
rect 69 387 75 393
rect 81 387 87 393
rect 93 387 99 393
rect 105 387 111 393
rect 117 387 123 393
rect 129 387 135 393
rect 141 387 147 393
rect 153 387 159 393
rect 165 387 171 393
rect 177 387 180 393
rect 0 384 180 387
rect 216 393 252 396
rect 216 387 219 393
rect 225 387 231 393
rect 237 387 243 393
rect 249 387 252 393
rect 216 384 252 387
rect 264 393 300 396
rect 264 387 267 393
rect 273 387 279 393
rect 285 387 291 393
rect 297 387 300 393
rect 264 384 300 387
rect 312 393 348 396
rect 312 387 315 393
rect 321 387 327 393
rect 333 387 339 393
rect 345 387 348 393
rect 312 384 348 387
rect 360 393 396 396
rect 360 387 363 393
rect 369 387 375 393
rect 381 387 387 393
rect 393 387 396 393
rect 360 384 396 387
rect 432 393 612 396
rect 432 387 435 393
rect 441 387 447 393
rect 453 387 459 393
rect 465 387 483 393
rect 489 387 495 393
rect 501 387 507 393
rect 513 387 519 393
rect 525 387 531 393
rect 537 387 543 393
rect 549 387 555 393
rect 561 387 579 393
rect 585 387 591 393
rect 597 387 603 393
rect 609 387 612 393
rect 432 384 612 387
rect 636 393 828 396
rect 636 387 639 393
rect 645 387 651 393
rect 657 387 663 393
rect 669 387 675 393
rect 681 387 699 393
rect 705 387 711 393
rect 717 387 723 393
rect 729 387 747 393
rect 753 387 759 393
rect 765 387 771 393
rect 777 387 795 393
rect 801 387 807 393
rect 813 387 819 393
rect 825 387 828 393
rect 636 384 828 387
rect 864 393 1044 396
rect 864 387 867 393
rect 873 387 879 393
rect 885 387 891 393
rect 897 387 903 393
rect 909 387 915 393
rect 921 387 927 393
rect 933 387 939 393
rect 945 387 963 393
rect 969 387 975 393
rect 981 387 987 393
rect 993 387 1011 393
rect 1017 387 1023 393
rect 1029 387 1035 393
rect 1041 387 1044 393
rect 864 384 1044 387
rect -12 357 0 360
rect -12 351 -9 357
rect -3 351 0 357
rect -12 345 0 351
rect -12 339 -9 345
rect -3 339 0 345
rect -12 333 0 339
rect -12 327 -9 333
rect -3 327 0 333
rect -12 324 0 327
rect 12 357 24 360
rect 12 351 15 357
rect 21 351 24 357
rect 12 345 24 351
rect 12 339 15 345
rect 21 339 24 345
rect 12 333 24 339
rect 12 327 15 333
rect 21 327 24 333
rect 12 324 24 327
rect 36 357 48 360
rect 36 351 39 357
rect 45 351 48 357
rect 36 345 48 351
rect 36 339 39 345
rect 45 339 48 345
rect 36 333 48 339
rect 36 327 39 333
rect 45 327 48 333
rect 36 324 48 327
rect 60 357 72 360
rect 60 351 63 357
rect 69 351 72 357
rect 60 345 72 351
rect 60 339 63 345
rect 69 339 72 345
rect 60 333 72 339
rect 60 327 63 333
rect 69 327 72 333
rect 60 324 72 327
rect 84 357 96 360
rect 84 351 87 357
rect 93 351 96 357
rect 84 345 96 351
rect 84 339 87 345
rect 93 339 96 345
rect 84 333 96 339
rect 84 327 87 333
rect 93 327 96 333
rect 84 324 96 327
rect 108 357 120 360
rect 108 351 111 357
rect 117 351 120 357
rect 108 345 120 351
rect 108 339 111 345
rect 117 339 120 345
rect 108 333 120 339
rect 108 327 111 333
rect 117 327 120 333
rect 108 324 120 327
rect 132 357 144 360
rect 132 351 135 357
rect 141 351 144 357
rect 132 345 144 351
rect 132 339 135 345
rect 141 339 144 345
rect 132 333 144 339
rect 132 327 135 333
rect 141 327 144 333
rect 132 324 144 327
rect 156 357 168 360
rect 156 351 159 357
rect 165 351 168 357
rect 156 345 168 351
rect 156 339 159 345
rect 165 339 168 345
rect 156 333 168 339
rect 156 327 159 333
rect 165 327 168 333
rect 156 324 168 327
rect 180 357 192 360
rect 180 351 183 357
rect 189 351 192 357
rect 180 345 192 351
rect 180 339 183 345
rect 189 339 192 345
rect 180 333 192 339
rect 180 327 183 333
rect 189 327 192 333
rect 180 324 192 327
rect 204 357 216 360
rect 204 351 207 357
rect 213 351 216 357
rect 204 345 216 351
rect 204 339 207 345
rect 213 339 216 345
rect 204 333 216 339
rect 204 327 207 333
rect 213 327 216 333
rect 204 324 216 327
rect 252 357 264 360
rect 252 351 255 357
rect 261 351 264 357
rect 252 345 264 351
rect 252 339 255 345
rect 261 339 264 345
rect 252 333 264 339
rect 252 327 255 333
rect 261 327 264 333
rect 252 324 264 327
rect 300 357 312 360
rect 300 351 303 357
rect 309 351 312 357
rect 300 345 312 351
rect 300 339 303 345
rect 309 339 312 345
rect 300 333 312 339
rect 300 327 303 333
rect 309 327 312 333
rect 300 324 312 327
rect 348 357 360 360
rect 348 351 351 357
rect 357 351 360 357
rect 348 345 360 351
rect 348 339 351 345
rect 357 339 360 345
rect 348 333 360 339
rect 348 327 351 333
rect 357 327 360 333
rect 348 324 360 327
rect 396 357 408 360
rect 396 351 399 357
rect 405 351 408 357
rect 396 345 408 351
rect 396 339 399 345
rect 405 339 408 345
rect 396 333 408 339
rect 396 327 399 333
rect 405 327 408 333
rect 396 324 408 327
rect 420 357 432 360
rect 420 351 423 357
rect 429 351 432 357
rect 420 345 432 351
rect 420 339 423 345
rect 429 339 432 345
rect 420 333 432 339
rect 420 327 423 333
rect 429 327 432 333
rect 420 324 432 327
rect 468 357 480 360
rect 468 351 471 357
rect 477 351 480 357
rect 468 345 480 351
rect 468 339 471 345
rect 477 339 480 345
rect 468 333 480 339
rect 468 327 471 333
rect 477 327 480 333
rect 468 324 480 327
rect 516 357 528 360
rect 516 351 519 357
rect 525 351 528 357
rect 516 345 528 351
rect 516 339 519 345
rect 525 339 528 345
rect 516 333 528 339
rect 516 327 519 333
rect 525 327 528 333
rect 516 324 528 327
rect 564 357 576 360
rect 564 351 567 357
rect 573 351 576 357
rect 564 345 576 351
rect 564 339 567 345
rect 573 339 576 345
rect 564 333 576 339
rect 564 327 567 333
rect 573 327 576 333
rect 564 324 576 327
rect 612 357 624 360
rect 612 351 615 357
rect 621 351 624 357
rect 612 345 624 351
rect 612 339 615 345
rect 621 339 624 345
rect 612 333 624 339
rect 612 327 615 333
rect 621 327 624 333
rect 612 324 624 327
rect 636 357 648 360
rect 636 351 639 357
rect 645 351 648 357
rect 636 345 648 351
rect 636 339 639 345
rect 645 339 648 345
rect 636 333 648 339
rect 636 327 639 333
rect 645 327 648 333
rect 636 324 648 327
rect 828 357 840 360
rect 828 351 831 357
rect 837 351 840 357
rect 828 345 840 351
rect 828 339 831 345
rect 837 339 840 345
rect 828 333 840 339
rect 828 327 831 333
rect 837 327 840 333
rect 828 324 840 327
rect 852 357 864 360
rect 852 351 855 357
rect 861 351 864 357
rect 852 345 864 351
rect 852 339 855 345
rect 861 339 864 345
rect 852 333 864 339
rect 852 327 855 333
rect 861 327 864 333
rect 852 324 864 327
rect 1044 357 1056 360
rect 1044 351 1047 357
rect 1053 351 1056 357
rect 1044 345 1056 351
rect 1044 339 1047 345
rect 1053 339 1056 345
rect 1044 333 1056 339
rect 1044 327 1047 333
rect 1053 327 1056 333
rect 1044 324 1056 327
rect 0 309 36 312
rect 0 303 3 309
rect 9 303 15 309
rect 21 303 27 309
rect 33 303 36 309
rect 0 300 36 303
rect 48 309 84 312
rect 48 303 51 309
rect 57 303 63 309
rect 69 303 75 309
rect 81 303 84 309
rect 48 300 84 303
rect 96 309 132 312
rect 96 303 99 309
rect 105 303 111 309
rect 117 303 123 309
rect 129 303 132 309
rect 96 300 132 303
rect 144 309 180 312
rect 144 303 147 309
rect 153 303 159 309
rect 165 303 171 309
rect 177 303 180 309
rect 144 300 180 303
rect 216 309 252 312
rect 216 303 219 309
rect 225 303 231 309
rect 237 303 243 309
rect 249 303 252 309
rect 216 300 252 303
rect 264 309 300 312
rect 264 303 267 309
rect 273 303 279 309
rect 285 303 291 309
rect 297 303 300 309
rect 264 300 300 303
rect 312 309 348 312
rect 312 303 315 309
rect 321 303 327 309
rect 333 303 339 309
rect 345 303 348 309
rect 312 300 348 303
rect 360 309 396 312
rect 360 303 363 309
rect 369 303 375 309
rect 381 303 387 309
rect 393 303 396 309
rect 360 300 396 303
rect 432 309 468 312
rect 432 303 435 309
rect 441 303 447 309
rect 453 303 459 309
rect 465 303 468 309
rect 432 300 468 303
rect 480 309 516 312
rect 480 303 483 309
rect 489 303 495 309
rect 501 303 507 309
rect 513 303 516 309
rect 480 300 516 303
rect 528 309 564 312
rect 528 303 531 309
rect 537 303 543 309
rect 549 303 555 309
rect 561 303 564 309
rect 528 300 564 303
rect 576 309 612 312
rect 576 303 579 309
rect 585 303 591 309
rect 597 303 603 309
rect 609 303 612 309
rect 576 300 612 303
rect 636 309 684 312
rect 636 303 639 309
rect 645 303 651 309
rect 657 303 663 309
rect 669 303 675 309
rect 681 303 684 309
rect 636 300 684 303
rect 696 309 732 312
rect 696 303 699 309
rect 705 303 711 309
rect 717 303 723 309
rect 729 303 732 309
rect 696 300 732 303
rect 744 309 780 312
rect 744 303 747 309
rect 753 303 759 309
rect 765 303 771 309
rect 777 303 780 309
rect 744 300 780 303
rect 792 309 840 312
rect 792 303 795 309
rect 801 303 807 309
rect 813 303 819 309
rect 825 303 831 309
rect 837 303 840 309
rect 792 300 840 303
rect 864 309 1044 312
rect 864 303 867 309
rect 873 303 879 309
rect 885 303 891 309
rect 897 303 903 309
rect 909 303 915 309
rect 921 303 927 309
rect 933 303 939 309
rect 945 303 963 309
rect 969 303 975 309
rect 981 303 987 309
rect 993 303 1011 309
rect 1017 303 1023 309
rect 1029 303 1035 309
rect 1041 303 1044 309
rect 864 300 1044 303
rect -12 285 1056 288
rect -12 279 -9 285
rect -3 279 3 285
rect 9 279 15 285
rect 21 279 27 285
rect 33 279 39 285
rect 45 279 51 285
rect 57 279 63 285
rect 69 279 75 285
rect 81 279 87 285
rect 93 279 99 285
rect 105 279 111 285
rect 117 279 123 285
rect 129 279 135 285
rect 141 279 147 285
rect 153 279 159 285
rect 165 279 171 285
rect 177 279 183 285
rect 189 279 195 285
rect 201 279 207 285
rect 213 279 219 285
rect 225 279 231 285
rect 237 279 243 285
rect 249 279 255 285
rect 261 279 267 285
rect 273 279 279 285
rect 285 279 291 285
rect 297 279 303 285
rect 309 279 315 285
rect 321 279 327 285
rect 333 279 339 285
rect 345 279 351 285
rect 357 279 363 285
rect 369 279 375 285
rect 381 279 387 285
rect 393 279 399 285
rect 405 279 411 285
rect 417 279 423 285
rect 429 279 435 285
rect 441 279 447 285
rect 453 279 459 285
rect 465 279 471 285
rect 477 279 483 285
rect 489 279 495 285
rect 501 279 507 285
rect 513 279 519 285
rect 525 279 531 285
rect 537 279 543 285
rect 549 279 555 285
rect 561 279 567 285
rect 573 279 579 285
rect 585 279 591 285
rect 597 279 603 285
rect 609 279 615 285
rect 621 279 627 285
rect 633 279 639 285
rect 645 279 651 285
rect 657 279 663 285
rect 669 279 675 285
rect 681 279 687 285
rect 693 279 699 285
rect 705 279 711 285
rect 717 279 723 285
rect 729 279 735 285
rect 741 279 747 285
rect 753 279 759 285
rect 765 279 771 285
rect 777 279 783 285
rect 789 279 795 285
rect 801 279 807 285
rect 813 279 819 285
rect 825 279 831 285
rect 837 279 843 285
rect 849 279 855 285
rect 861 279 867 285
rect 873 279 879 285
rect 885 279 891 285
rect 897 279 903 285
rect 909 279 915 285
rect 921 279 927 285
rect 933 279 939 285
rect 945 279 951 285
rect 957 279 963 285
rect 969 279 975 285
rect 981 279 987 285
rect 993 279 999 285
rect 1005 279 1011 285
rect 1017 279 1023 285
rect 1029 279 1035 285
rect 1041 279 1047 285
rect 1053 279 1056 285
rect -12 276 1056 279
rect -24 261 1056 264
rect -24 255 -21 261
rect -15 255 -9 261
rect -3 255 3 261
rect 9 255 15 261
rect 21 255 27 261
rect 33 255 39 261
rect 45 255 51 261
rect 57 255 63 261
rect 69 255 75 261
rect 81 255 87 261
rect 93 255 99 261
rect 105 255 111 261
rect 117 255 123 261
rect 129 255 135 261
rect 141 255 147 261
rect 153 255 159 261
rect 165 255 171 261
rect 177 255 183 261
rect 189 255 195 261
rect 201 255 207 261
rect 213 255 219 261
rect 225 255 231 261
rect 237 255 243 261
rect 249 255 255 261
rect 261 255 267 261
rect 273 255 279 261
rect 285 255 291 261
rect 297 255 303 261
rect 309 255 315 261
rect 321 255 327 261
rect 333 255 339 261
rect 345 255 351 261
rect 357 255 363 261
rect 369 255 375 261
rect 381 255 387 261
rect 393 255 399 261
rect 405 255 411 261
rect 417 255 423 261
rect 429 255 435 261
rect 441 255 447 261
rect 453 255 459 261
rect 465 255 471 261
rect 477 255 483 261
rect 489 255 495 261
rect 501 255 507 261
rect 513 255 519 261
rect 525 255 531 261
rect 537 255 543 261
rect 549 255 555 261
rect 561 255 567 261
rect 573 255 579 261
rect 585 255 591 261
rect 597 255 603 261
rect 609 255 615 261
rect 621 255 627 261
rect 633 255 639 261
rect 645 255 651 261
rect 657 255 663 261
rect 669 255 675 261
rect 681 255 687 261
rect 693 255 699 261
rect 705 255 711 261
rect 717 255 723 261
rect 729 255 735 261
rect 741 255 747 261
rect 753 255 759 261
rect 765 255 771 261
rect 777 255 783 261
rect 789 255 795 261
rect 801 255 807 261
rect 813 255 819 261
rect 825 255 831 261
rect 837 255 843 261
rect 849 255 855 261
rect 861 255 867 261
rect 873 255 879 261
rect 885 255 891 261
rect 897 255 903 261
rect 909 255 915 261
rect 921 255 927 261
rect 933 255 939 261
rect 945 255 951 261
rect 957 255 963 261
rect 969 255 975 261
rect 981 255 987 261
rect 993 255 999 261
rect 1005 255 1011 261
rect 1017 255 1023 261
rect 1029 255 1035 261
rect 1041 255 1047 261
rect 1053 255 1056 261
rect -24 252 1056 255
rect -12 237 192 240
rect -12 231 -9 237
rect -3 231 3 237
rect 9 231 15 237
rect 21 231 27 237
rect 33 231 39 237
rect 45 231 51 237
rect 57 231 63 237
rect 69 231 75 237
rect 81 231 87 237
rect 93 231 99 237
rect 105 231 111 237
rect 117 231 123 237
rect 129 231 135 237
rect 141 231 147 237
rect 153 231 159 237
rect 165 231 171 237
rect 177 231 183 237
rect 189 231 192 237
rect -12 228 192 231
rect 216 237 252 240
rect 216 231 219 237
rect 225 231 231 237
rect 237 231 243 237
rect 249 231 252 237
rect 216 228 252 231
rect 264 237 300 240
rect 264 231 267 237
rect 273 231 279 237
rect 285 231 291 237
rect 297 231 300 237
rect 264 228 300 231
rect 312 237 348 240
rect 312 231 315 237
rect 321 231 327 237
rect 333 231 339 237
rect 345 231 348 237
rect 312 228 348 231
rect 360 237 396 240
rect 360 231 363 237
rect 369 231 375 237
rect 381 231 387 237
rect 393 231 396 237
rect 360 228 396 231
rect 432 237 468 240
rect 432 231 435 237
rect 441 231 447 237
rect 453 231 459 237
rect 465 231 468 237
rect 432 228 468 231
rect 480 237 516 240
rect 480 231 483 237
rect 489 231 495 237
rect 501 231 507 237
rect 513 231 516 237
rect 480 228 516 231
rect 528 237 564 240
rect 528 231 531 237
rect 537 231 543 237
rect 549 231 555 237
rect 561 231 564 237
rect 528 228 564 231
rect 576 237 612 240
rect 576 231 579 237
rect 585 231 591 237
rect 597 231 603 237
rect 609 231 612 237
rect 576 228 612 231
rect 648 237 684 240
rect 648 231 651 237
rect 657 231 663 237
rect 669 231 675 237
rect 681 231 684 237
rect 648 228 684 231
rect 696 237 732 240
rect 696 231 699 237
rect 705 231 711 237
rect 717 231 723 237
rect 729 231 732 237
rect 696 228 732 231
rect 744 237 780 240
rect 744 231 747 237
rect 753 231 759 237
rect 765 231 771 237
rect 777 231 780 237
rect 744 228 780 231
rect 792 237 828 240
rect 792 231 795 237
rect 801 231 807 237
rect 813 231 819 237
rect 825 231 828 237
rect 792 228 828 231
rect 864 237 876 240
rect 864 231 867 237
rect 873 231 876 237
rect 864 228 876 231
rect 912 237 948 240
rect 912 231 915 237
rect 921 231 927 237
rect 933 231 939 237
rect 945 231 948 237
rect 912 228 948 231
rect 960 237 996 240
rect 960 231 963 237
rect 969 231 975 237
rect 981 231 987 237
rect 993 231 996 237
rect 960 228 996 231
rect 1008 237 1044 240
rect 1008 231 1011 237
rect 1017 231 1023 237
rect 1029 231 1035 237
rect 1041 231 1044 237
rect 1008 228 1044 231
rect 1080 237 1116 240
rect 1080 231 1083 237
rect 1089 231 1095 237
rect 1101 231 1107 237
rect 1113 231 1116 237
rect 1080 228 1116 231
rect 1128 237 1164 240
rect 1128 231 1131 237
rect 1137 231 1143 237
rect 1149 231 1155 237
rect 1161 231 1164 237
rect 1128 228 1164 231
rect 1176 237 1212 240
rect 1176 231 1179 237
rect 1185 231 1191 237
rect 1197 231 1203 237
rect 1209 231 1212 237
rect 1176 228 1212 231
rect 1224 237 1260 240
rect 1224 231 1227 237
rect 1233 231 1239 237
rect 1245 231 1251 237
rect 1257 231 1260 237
rect 1224 228 1260 231
rect -12 213 0 216
rect -12 207 -9 213
rect -3 207 0 213
rect -12 201 0 207
rect -12 195 -9 201
rect -3 195 0 201
rect -12 189 0 195
rect -12 183 -9 189
rect -3 183 0 189
rect -12 180 0 183
rect 12 213 24 228
rect 12 207 15 213
rect 21 207 24 213
rect 12 201 24 207
rect 12 195 15 201
rect 21 195 24 201
rect 12 189 24 195
rect 12 183 15 189
rect 21 183 24 189
rect 12 180 24 183
rect 36 213 48 216
rect 36 207 39 213
rect 45 207 48 213
rect 36 201 48 207
rect 36 195 39 201
rect 45 195 48 201
rect 36 189 48 195
rect 36 183 39 189
rect 45 183 48 189
rect 36 180 48 183
rect 60 213 72 228
rect 60 207 63 213
rect 69 207 72 213
rect 60 201 72 207
rect 60 195 63 201
rect 69 195 72 201
rect 60 189 72 195
rect 60 183 63 189
rect 69 183 72 189
rect 60 180 72 183
rect 84 213 96 216
rect 84 207 87 213
rect 93 207 96 213
rect 84 201 96 207
rect 84 195 87 201
rect 93 195 96 201
rect 84 189 96 195
rect 84 183 87 189
rect 93 183 96 189
rect 84 180 96 183
rect 108 213 120 228
rect 108 207 111 213
rect 117 207 120 213
rect 108 201 120 207
rect 108 195 111 201
rect 117 195 120 201
rect 108 189 120 195
rect 108 183 111 189
rect 117 183 120 189
rect 108 180 120 183
rect 132 213 144 216
rect 132 207 135 213
rect 141 207 144 213
rect 132 201 144 207
rect 132 195 135 201
rect 141 195 144 201
rect 132 189 144 195
rect 132 183 135 189
rect 141 183 144 189
rect 132 180 144 183
rect 156 213 168 228
rect 156 207 159 213
rect 165 207 168 213
rect 156 201 168 207
rect 156 195 159 201
rect 165 195 168 201
rect 156 189 168 195
rect 156 183 159 189
rect 165 183 168 189
rect 156 180 168 183
rect 180 213 192 216
rect 180 207 183 213
rect 189 207 192 213
rect 180 201 192 207
rect 180 195 183 201
rect 189 195 192 201
rect 180 189 192 195
rect 180 183 183 189
rect 189 183 192 189
rect 180 180 192 183
rect 204 213 216 216
rect 204 207 207 213
rect 213 207 216 213
rect 204 201 216 207
rect 204 195 207 201
rect 213 195 216 201
rect 204 189 216 195
rect 204 183 207 189
rect 213 183 216 189
rect 204 180 216 183
rect 300 213 312 216
rect 300 207 303 213
rect 309 207 312 213
rect 300 201 312 207
rect 300 195 303 201
rect 309 195 312 201
rect 300 189 312 195
rect 300 183 303 189
rect 309 183 312 189
rect 300 180 312 183
rect 396 213 408 216
rect 396 207 399 213
rect 405 207 408 213
rect 396 201 408 207
rect 396 195 399 201
rect 405 195 408 201
rect 396 189 408 195
rect 396 183 399 189
rect 405 183 408 189
rect 396 180 408 183
rect 420 213 432 216
rect 420 207 423 213
rect 429 207 432 213
rect 420 201 432 207
rect 420 195 423 201
rect 429 195 432 201
rect 420 189 432 195
rect 420 183 423 189
rect 429 183 432 189
rect 420 180 432 183
rect 516 213 528 216
rect 516 207 519 213
rect 525 207 528 213
rect 516 201 528 207
rect 516 195 519 201
rect 525 195 528 201
rect 516 189 528 195
rect 516 183 519 189
rect 525 183 528 189
rect 516 180 528 183
rect 612 213 624 216
rect 612 207 615 213
rect 621 207 624 213
rect 612 201 624 207
rect 612 195 615 201
rect 621 195 624 201
rect 612 189 624 195
rect 612 183 615 189
rect 621 183 624 189
rect 612 180 624 183
rect 636 213 648 216
rect 636 207 639 213
rect 645 207 648 213
rect 636 201 648 207
rect 636 195 639 201
rect 645 195 648 201
rect 636 189 648 195
rect 636 183 639 189
rect 645 183 648 189
rect 636 180 648 183
rect 732 213 744 216
rect 732 207 735 213
rect 741 207 744 213
rect 732 201 744 207
rect 732 195 735 201
rect 741 195 744 201
rect 732 189 744 195
rect 732 183 735 189
rect 741 183 744 189
rect 732 180 744 183
rect 828 213 840 216
rect 828 207 831 213
rect 837 207 840 213
rect 828 201 840 207
rect 828 195 831 201
rect 837 195 840 201
rect 828 189 840 195
rect 828 183 831 189
rect 837 183 840 189
rect 828 180 840 183
rect 852 213 864 216
rect 852 207 855 213
rect 861 207 864 213
rect 852 201 864 207
rect 852 195 855 201
rect 861 195 864 201
rect 852 189 864 195
rect 852 183 855 189
rect 861 183 864 189
rect 852 180 864 183
rect 876 213 888 216
rect 876 207 879 213
rect 885 207 888 213
rect 876 201 888 207
rect 876 195 879 201
rect 885 195 888 201
rect 876 189 888 195
rect 876 183 879 189
rect 885 183 888 189
rect 876 180 888 183
rect 900 213 912 216
rect 900 207 903 213
rect 909 207 912 213
rect 900 201 912 207
rect 900 195 903 201
rect 909 195 912 201
rect 900 189 912 195
rect 900 183 903 189
rect 909 183 912 189
rect 900 180 912 183
rect 1044 213 1056 216
rect 1044 207 1047 213
rect 1053 207 1056 213
rect 1044 201 1056 207
rect 1044 195 1047 201
rect 1053 195 1056 201
rect 1044 189 1056 195
rect 1044 183 1047 189
rect 1053 183 1056 189
rect 1044 180 1056 183
rect 1068 213 1080 216
rect 1068 207 1071 213
rect 1077 207 1080 213
rect 1068 201 1080 207
rect 1068 195 1071 201
rect 1077 195 1080 201
rect 1068 189 1080 195
rect 1068 183 1071 189
rect 1077 183 1080 189
rect 1068 180 1080 183
rect 1164 213 1176 216
rect 1164 207 1167 213
rect 1173 207 1176 213
rect 1164 201 1176 207
rect 1164 195 1167 201
rect 1173 195 1176 201
rect 1164 189 1176 195
rect 1164 183 1167 189
rect 1173 183 1176 189
rect 1164 180 1176 183
rect 1260 213 1272 216
rect 1260 207 1263 213
rect 1269 207 1272 213
rect 1260 201 1272 207
rect 1260 195 1263 201
rect 1269 195 1272 201
rect 1260 189 1272 195
rect 1260 183 1263 189
rect 1269 183 1272 189
rect 1260 180 1272 183
rect 0 69 36 72
rect 0 63 3 69
rect 9 63 15 69
rect 21 63 27 69
rect 33 63 36 69
rect 0 60 36 63
rect 48 69 84 72
rect 48 63 51 69
rect 57 63 63 69
rect 69 63 75 69
rect 81 63 84 69
rect 48 60 84 63
rect 96 69 132 72
rect 96 63 99 69
rect 105 63 111 69
rect 117 63 123 69
rect 129 63 132 69
rect 96 60 132 63
rect 144 69 180 72
rect 144 63 147 69
rect 153 63 159 69
rect 165 63 171 69
rect 177 63 180 69
rect 144 60 180 63
rect 216 69 252 72
rect 216 63 219 69
rect 225 63 231 69
rect 237 63 243 69
rect 249 63 252 69
rect 216 60 252 63
rect 264 69 300 72
rect 264 63 267 69
rect 273 63 279 69
rect 285 63 291 69
rect 297 63 300 69
rect 264 60 300 63
rect 312 69 348 72
rect 312 63 315 69
rect 321 63 327 69
rect 333 63 339 69
rect 345 63 348 69
rect 312 60 348 63
rect 360 69 396 72
rect 360 63 363 69
rect 369 63 375 69
rect 381 63 387 69
rect 393 63 396 69
rect 360 60 396 63
rect 432 69 468 72
rect 432 63 435 69
rect 441 63 447 69
rect 453 63 459 69
rect 465 63 468 69
rect 432 60 468 63
rect 480 69 516 72
rect 480 63 483 69
rect 489 63 495 69
rect 501 63 507 69
rect 513 63 516 69
rect 480 60 516 63
rect 528 69 564 72
rect 528 63 531 69
rect 537 63 543 69
rect 549 63 555 69
rect 561 63 564 69
rect 528 60 564 63
rect 576 69 612 72
rect 576 63 579 69
rect 585 63 591 69
rect 597 63 603 69
rect 609 63 612 69
rect 576 60 612 63
rect 648 69 684 72
rect 648 63 651 69
rect 657 63 663 69
rect 669 63 675 69
rect 681 63 684 69
rect 648 60 684 63
rect 696 69 732 72
rect 696 63 699 69
rect 705 63 711 69
rect 717 63 723 69
rect 729 63 732 69
rect 696 60 732 63
rect 744 69 780 72
rect 744 63 747 69
rect 753 63 759 69
rect 765 63 771 69
rect 777 63 780 69
rect 744 60 780 63
rect 792 69 828 72
rect 792 63 795 69
rect 801 63 807 69
rect 813 63 819 69
rect 825 63 828 69
rect 792 60 828 63
rect 864 69 900 72
rect 864 63 867 69
rect 873 63 879 69
rect 885 63 891 69
rect 897 63 900 69
rect 864 60 900 63
rect 912 69 948 72
rect 912 63 915 69
rect 921 63 927 69
rect 933 63 939 69
rect 945 63 948 69
rect 912 60 948 63
rect 960 69 996 72
rect 960 63 963 69
rect 969 63 975 69
rect 981 63 987 69
rect 993 63 996 69
rect 960 60 996 63
rect 1008 69 1044 72
rect 1008 63 1011 69
rect 1017 63 1023 69
rect 1029 63 1035 69
rect 1041 63 1044 69
rect 1008 60 1044 63
rect 1080 69 1116 72
rect 1080 63 1083 69
rect 1089 63 1095 69
rect 1101 63 1107 69
rect 1113 63 1116 69
rect 1080 60 1116 63
rect 1128 69 1164 72
rect 1128 63 1131 69
rect 1137 63 1143 69
rect 1149 63 1155 69
rect 1161 63 1164 69
rect 1128 60 1164 63
rect 1176 69 1212 72
rect 1176 63 1179 69
rect 1185 63 1191 69
rect 1197 63 1203 69
rect 1209 63 1212 69
rect 1176 60 1212 63
rect 1224 69 1260 72
rect 1224 63 1227 69
rect 1233 63 1239 69
rect 1245 63 1251 69
rect 1257 63 1260 69
rect 1224 60 1260 63
rect -12 45 0 48
rect -12 39 -9 45
rect -3 39 0 45
rect -12 33 0 39
rect -12 27 -9 33
rect -3 27 0 33
rect -12 21 0 27
rect -12 15 -9 21
rect -3 15 0 21
rect -12 0 0 15
rect 36 45 48 48
rect 36 39 39 45
rect 45 39 48 45
rect 36 33 48 39
rect 36 27 39 33
rect 45 27 48 33
rect 36 21 48 27
rect 36 15 39 21
rect 45 15 48 21
rect 36 12 48 15
rect 84 45 96 48
rect 84 39 87 45
rect 93 39 96 45
rect 84 33 96 39
rect 84 27 87 33
rect 93 27 96 33
rect 84 21 96 27
rect 84 15 87 21
rect 93 15 96 21
rect 84 12 96 15
rect 132 45 144 48
rect 132 39 135 45
rect 141 39 144 45
rect 132 33 144 39
rect 132 27 135 33
rect 141 27 144 33
rect 132 21 144 27
rect 132 15 135 21
rect 141 15 144 21
rect 132 12 144 15
rect 180 45 192 48
rect 180 39 183 45
rect 189 39 192 45
rect 180 33 192 39
rect 180 27 183 33
rect 189 27 192 33
rect 180 21 192 27
rect 180 15 183 21
rect 189 15 192 21
rect 180 0 192 15
rect 204 45 216 48
rect 204 39 207 45
rect 213 39 216 45
rect 204 33 216 39
rect 204 27 207 33
rect 213 27 216 33
rect 204 21 216 27
rect 204 15 207 21
rect 213 15 216 21
rect 204 0 216 15
rect 252 45 264 48
rect 252 39 255 45
rect 261 39 264 45
rect 252 33 264 39
rect 252 27 255 33
rect 261 27 264 33
rect 252 21 264 27
rect 252 15 255 21
rect 261 15 264 21
rect 252 12 264 15
rect 300 45 312 48
rect 300 39 303 45
rect 309 39 312 45
rect 300 33 312 39
rect 300 27 303 33
rect 309 27 312 33
rect 300 21 312 27
rect 300 15 303 21
rect 309 15 312 21
rect 300 12 312 15
rect 348 45 360 48
rect 348 39 351 45
rect 357 39 360 45
rect 348 33 360 39
rect 348 27 351 33
rect 357 27 360 33
rect 348 21 360 27
rect 348 15 351 21
rect 357 15 360 21
rect 348 12 360 15
rect 396 45 408 48
rect 396 39 399 45
rect 405 39 408 45
rect 396 33 408 39
rect 396 27 399 33
rect 405 27 408 33
rect 396 21 408 27
rect 396 15 399 21
rect 405 15 408 21
rect 396 0 408 15
rect 420 45 432 48
rect 420 39 423 45
rect 429 39 432 45
rect 420 33 432 39
rect 420 27 423 33
rect 429 27 432 33
rect 420 21 432 27
rect 420 15 423 21
rect 429 15 432 21
rect 420 0 432 15
rect 516 45 528 48
rect 516 39 519 45
rect 525 39 528 45
rect 516 33 528 39
rect 516 27 519 33
rect 525 27 528 33
rect 516 21 528 27
rect 516 15 519 21
rect 525 15 528 21
rect 516 12 528 15
rect 612 45 624 48
rect 612 39 615 45
rect 621 39 624 45
rect 612 33 624 39
rect 612 27 615 33
rect 621 27 624 33
rect 612 21 624 27
rect 612 15 615 21
rect 621 15 624 21
rect 612 0 624 15
rect 636 45 648 48
rect 636 39 639 45
rect 645 39 648 45
rect 636 33 648 39
rect 636 27 639 33
rect 645 27 648 33
rect 636 21 648 27
rect 636 15 639 21
rect 645 15 648 21
rect 636 0 648 15
rect 732 45 744 48
rect 732 39 735 45
rect 741 39 744 45
rect 732 33 744 39
rect 732 27 735 33
rect 741 27 744 33
rect 732 21 744 27
rect 732 15 735 21
rect 741 15 744 21
rect 732 12 744 15
rect 828 45 840 48
rect 828 39 831 45
rect 837 39 840 45
rect 828 33 840 39
rect 828 27 831 33
rect 837 27 840 33
rect 828 21 840 27
rect 828 15 831 21
rect 837 15 840 21
rect 828 0 840 15
rect 852 45 864 48
rect 852 39 855 45
rect 861 39 864 45
rect 852 33 864 39
rect 852 27 855 33
rect 861 27 864 33
rect 852 21 864 27
rect 852 15 855 21
rect 861 15 864 21
rect 852 0 864 15
rect 1044 45 1056 48
rect 1044 39 1047 45
rect 1053 39 1056 45
rect 1044 33 1056 39
rect 1044 27 1047 33
rect 1053 27 1056 33
rect 1044 21 1056 27
rect 1044 15 1047 21
rect 1053 15 1056 21
rect 1044 12 1056 15
rect 1068 45 1080 48
rect 1068 39 1071 45
rect 1077 39 1080 45
rect 1068 33 1080 39
rect 1068 27 1071 33
rect 1077 27 1080 33
rect 1068 21 1080 27
rect 1068 15 1071 21
rect 1077 15 1080 21
rect 1068 0 1080 15
rect 1164 45 1176 48
rect 1164 39 1167 45
rect 1173 39 1176 45
rect 1164 33 1176 39
rect 1164 27 1167 33
rect 1173 27 1176 33
rect 1164 21 1176 27
rect 1164 15 1167 21
rect 1173 15 1176 21
rect 1164 12 1176 15
rect 1260 45 1272 48
rect 1260 39 1263 45
rect 1269 39 1272 45
rect 1260 33 1272 39
rect 1260 27 1263 33
rect 1269 27 1272 33
rect 1260 21 1272 27
rect 1260 15 1263 21
rect 1269 15 1272 21
rect 1260 0 1272 15
rect -24 -3 1272 0
rect -24 -9 -21 -3
rect -15 -9 -9 -3
rect -3 -9 3 -3
rect 9 -9 15 -3
rect 21 -9 27 -3
rect 33 -9 39 -3
rect 45 -9 51 -3
rect 57 -9 63 -3
rect 69 -9 75 -3
rect 81 -9 87 -3
rect 93 -9 99 -3
rect 105 -9 111 -3
rect 117 -9 123 -3
rect 129 -9 135 -3
rect 141 -9 147 -3
rect 153 -9 159 -3
rect 165 -9 171 -3
rect 177 -9 183 -3
rect 189 -9 195 -3
rect 201 -9 207 -3
rect 213 -9 219 -3
rect 225 -9 231 -3
rect 237 -9 243 -3
rect 249 -9 255 -3
rect 261 -9 267 -3
rect 273 -9 279 -3
rect 285 -9 291 -3
rect 297 -9 303 -3
rect 309 -9 315 -3
rect 321 -9 327 -3
rect 333 -9 339 -3
rect 345 -9 351 -3
rect 357 -9 363 -3
rect 369 -9 375 -3
rect 381 -9 387 -3
rect 393 -9 399 -3
rect 405 -9 411 -3
rect 417 -9 423 -3
rect 429 -9 435 -3
rect 441 -9 447 -3
rect 453 -9 459 -3
rect 465 -9 471 -3
rect 477 -9 483 -3
rect 489 -9 495 -3
rect 501 -9 507 -3
rect 513 -9 519 -3
rect 525 -9 531 -3
rect 537 -9 543 -3
rect 549 -9 555 -3
rect 561 -9 567 -3
rect 573 -9 579 -3
rect 585 -9 591 -3
rect 597 -9 603 -3
rect 609 -9 615 -3
rect 621 -9 627 -3
rect 633 -9 639 -3
rect 645 -9 651 -3
rect 657 -9 663 -3
rect 669 -9 675 -3
rect 681 -9 687 -3
rect 693 -9 699 -3
rect 705 -9 711 -3
rect 717 -9 723 -3
rect 729 -9 735 -3
rect 741 -9 747 -3
rect 753 -9 759 -3
rect 765 -9 771 -3
rect 777 -9 783 -3
rect 789 -9 795 -3
rect 801 -9 807 -3
rect 813 -9 819 -3
rect 825 -9 831 -3
rect 837 -9 843 -3
rect 849 -9 855 -3
rect 861 -9 867 -3
rect 873 -9 879 -3
rect 885 -9 891 -3
rect 897 -9 903 -3
rect 909 -9 915 -3
rect 921 -9 927 -3
rect 933 -9 939 -3
rect 945 -9 951 -3
rect 957 -9 963 -3
rect 969 -9 975 -3
rect 981 -9 987 -3
rect 993 -9 999 -3
rect 1005 -9 1011 -3
rect 1017 -9 1023 -3
rect 1029 -9 1035 -3
rect 1041 -9 1047 -3
rect 1053 -9 1059 -3
rect 1065 -9 1071 -3
rect 1077 -9 1083 -3
rect 1089 -9 1095 -3
rect 1101 -9 1107 -3
rect 1113 -9 1119 -3
rect 1125 -9 1131 -3
rect 1137 -9 1143 -3
rect 1149 -9 1155 -3
rect 1161 -9 1167 -3
rect 1173 -9 1179 -3
rect 1185 -9 1191 -3
rect 1197 -9 1203 -3
rect 1209 -9 1215 -3
rect 1221 -9 1227 -3
rect 1233 -9 1239 -3
rect 1245 -9 1251 -3
rect 1257 -9 1263 -3
rect 1269 -9 1272 -3
rect -24 -12 1272 -9
<< via1 >>
rect -9 435 -3 441
rect -9 423 -3 429
rect -9 411 -3 417
rect 15 435 21 441
rect 15 423 21 429
rect 15 411 21 417
rect 39 435 45 441
rect 39 423 45 429
rect 39 411 45 417
rect 63 435 69 441
rect 63 423 69 429
rect 63 411 69 417
rect 87 435 93 441
rect 87 423 93 429
rect 87 411 93 417
rect 111 435 117 441
rect 111 423 117 429
rect 111 411 117 417
rect 135 435 141 441
rect 135 423 141 429
rect 135 411 141 417
rect 159 435 165 441
rect 159 423 165 429
rect 159 411 165 417
rect 183 435 189 441
rect 183 423 189 429
rect 183 411 189 417
rect 207 435 213 441
rect 207 423 213 429
rect 207 411 213 417
rect 255 435 261 441
rect 255 423 261 429
rect 255 411 261 417
rect 303 435 309 441
rect 303 423 309 429
rect 303 411 309 417
rect 351 435 357 441
rect 351 423 357 429
rect 351 411 357 417
rect 399 435 405 441
rect 399 423 405 429
rect 399 411 405 417
rect 423 435 429 441
rect 423 423 429 429
rect 423 411 429 417
rect 471 435 477 441
rect 471 423 477 429
rect 471 411 477 417
rect 519 435 525 441
rect 519 423 525 429
rect 519 411 525 417
rect 567 435 573 441
rect 567 423 573 429
rect 567 411 573 417
rect 615 435 621 441
rect 615 423 621 429
rect 615 411 621 417
rect 639 435 645 441
rect 639 423 645 429
rect 639 411 645 417
rect 831 435 837 441
rect 831 423 837 429
rect 831 411 837 417
rect 855 435 861 441
rect 855 423 861 429
rect 855 411 861 417
rect 1047 435 1053 441
rect 1047 423 1053 429
rect 1047 411 1053 417
rect 39 387 45 393
rect 87 387 93 393
rect 135 387 141 393
rect 231 387 237 393
rect 279 387 285 393
rect 327 387 333 393
rect 375 387 381 393
rect 519 387 525 393
rect 639 387 645 393
rect 903 387 909 393
rect -9 351 -3 357
rect -9 339 -3 345
rect -9 327 -3 333
rect 15 351 21 357
rect 15 339 21 345
rect 15 327 21 333
rect 39 351 45 357
rect 39 339 45 345
rect 39 327 45 333
rect 63 351 69 357
rect 63 339 69 345
rect 63 327 69 333
rect 87 351 93 357
rect 87 339 93 345
rect 87 327 93 333
rect 111 351 117 357
rect 111 339 117 345
rect 111 327 117 333
rect 135 351 141 357
rect 135 339 141 345
rect 135 327 141 333
rect 159 351 165 357
rect 159 339 165 345
rect 159 327 165 333
rect 183 351 189 357
rect 183 339 189 345
rect 183 327 189 333
rect 207 351 213 357
rect 207 339 213 345
rect 207 327 213 333
rect 255 351 261 357
rect 255 339 261 345
rect 255 327 261 333
rect 303 351 309 357
rect 303 339 309 345
rect 303 327 309 333
rect 351 351 357 357
rect 351 339 357 345
rect 351 327 357 333
rect 399 351 405 357
rect 399 339 405 345
rect 399 327 405 333
rect 423 351 429 357
rect 423 339 429 345
rect 423 327 429 333
rect 471 351 477 357
rect 471 339 477 345
rect 471 327 477 333
rect 519 351 525 357
rect 519 339 525 345
rect 519 327 525 333
rect 567 351 573 357
rect 567 339 573 345
rect 567 327 573 333
rect 615 351 621 357
rect 615 339 621 345
rect 615 327 621 333
rect 639 351 645 357
rect 639 339 645 345
rect 639 327 645 333
rect 831 351 837 357
rect 831 339 837 345
rect 831 327 837 333
rect 855 351 861 357
rect 855 339 861 345
rect 855 327 861 333
rect 1047 351 1053 357
rect 1047 339 1053 345
rect 1047 327 1053 333
rect 15 303 21 309
rect 63 303 69 309
rect 111 303 117 309
rect 159 303 165 309
rect 231 303 237 309
rect 279 303 285 309
rect 327 303 333 309
rect 375 303 381 309
rect 447 303 453 309
rect 495 303 501 309
rect 543 303 549 309
rect 591 303 597 309
rect 639 303 645 309
rect 663 303 669 309
rect 711 303 717 309
rect 759 303 765 309
rect 807 303 813 309
rect 831 303 837 309
rect 903 303 909 309
rect -9 231 -3 237
rect 39 231 45 237
rect 87 231 93 237
rect 135 231 141 237
rect 183 231 189 237
rect 231 231 237 237
rect 279 231 285 237
rect 327 231 333 237
rect 375 231 381 237
rect 447 231 453 237
rect 495 231 501 237
rect 543 231 549 237
rect 591 231 597 237
rect 663 231 669 237
rect 711 231 717 237
rect 759 231 765 237
rect 807 231 813 237
rect 867 231 873 237
rect 927 231 933 237
rect 975 231 981 237
rect 1023 231 1029 237
rect 1095 231 1101 237
rect 1143 231 1149 237
rect 1191 231 1197 237
rect 1239 231 1245 237
rect -9 207 -3 213
rect -9 195 -3 201
rect -9 183 -3 189
rect 39 207 45 213
rect 39 195 45 201
rect 39 183 45 189
rect 87 207 93 213
rect 87 195 93 201
rect 87 183 93 189
rect 135 207 141 213
rect 135 195 141 201
rect 135 183 141 189
rect 183 207 189 213
rect 183 195 189 201
rect 183 183 189 189
rect 207 207 213 213
rect 207 195 213 201
rect 207 183 213 189
rect 303 207 309 213
rect 303 195 309 201
rect 303 183 309 189
rect 399 207 405 213
rect 399 195 405 201
rect 399 183 405 189
rect 423 207 429 213
rect 423 195 429 201
rect 423 183 429 189
rect 519 207 525 213
rect 519 195 525 201
rect 519 183 525 189
rect 615 207 621 213
rect 615 195 621 201
rect 615 183 621 189
rect 639 207 645 213
rect 639 195 645 201
rect 639 183 645 189
rect 735 207 741 213
rect 735 195 741 201
rect 735 183 741 189
rect 831 207 837 213
rect 831 195 837 201
rect 831 183 837 189
rect 855 207 861 213
rect 855 195 861 201
rect 855 183 861 189
rect 879 207 885 213
rect 879 195 885 201
rect 879 183 885 189
rect 903 207 909 213
rect 903 195 909 201
rect 903 183 909 189
rect 1047 207 1053 213
rect 1047 195 1053 201
rect 1047 183 1053 189
rect 1071 207 1077 213
rect 1071 195 1077 201
rect 1071 183 1077 189
rect 1167 207 1173 213
rect 1167 195 1173 201
rect 1167 183 1173 189
rect 1263 207 1269 213
rect 1263 195 1269 201
rect 1263 183 1269 189
rect 15 63 21 69
rect 63 63 69 69
rect 111 63 117 69
rect 159 63 165 69
rect 231 63 237 69
rect 279 63 285 69
rect 327 63 333 69
rect 375 63 381 69
rect 447 63 453 69
rect 495 63 501 69
rect 543 63 549 69
rect 591 63 597 69
rect 663 63 669 69
rect 711 63 717 69
rect 759 63 765 69
rect 807 63 813 69
rect 879 63 885 69
rect 927 63 933 69
rect 975 63 981 69
rect 1023 63 1029 69
rect 1095 63 1101 69
rect 1143 63 1149 69
rect 1191 63 1197 69
rect 1239 63 1245 69
rect -9 39 -3 45
rect -9 27 -3 33
rect -9 15 -3 21
rect 39 39 45 45
rect 39 27 45 33
rect 39 15 45 21
rect 87 39 93 45
rect 87 27 93 33
rect 87 15 93 21
rect 135 39 141 45
rect 135 27 141 33
rect 135 15 141 21
rect 183 39 189 45
rect 183 27 189 33
rect 183 15 189 21
rect 207 39 213 45
rect 207 27 213 33
rect 207 15 213 21
rect 255 39 261 45
rect 255 27 261 33
rect 255 15 261 21
rect 303 39 309 45
rect 303 27 309 33
rect 303 15 309 21
rect 351 39 357 45
rect 351 27 357 33
rect 351 15 357 21
rect 399 39 405 45
rect 399 27 405 33
rect 399 15 405 21
rect 423 39 429 45
rect 423 27 429 33
rect 423 15 429 21
rect 519 39 525 45
rect 519 27 525 33
rect 519 15 525 21
rect 615 39 621 45
rect 615 27 621 33
rect 615 15 621 21
rect 639 39 645 45
rect 639 27 645 33
rect 639 15 645 21
rect 735 39 741 45
rect 735 27 741 33
rect 735 15 741 21
rect 831 39 837 45
rect 831 27 837 33
rect 831 15 837 21
rect 855 39 861 45
rect 855 27 861 33
rect 855 15 861 21
rect 1047 39 1053 45
rect 1047 27 1053 33
rect 1047 15 1053 21
rect 1071 39 1077 45
rect 1071 27 1077 33
rect 1071 15 1077 21
rect 1167 39 1173 45
rect 1167 27 1173 33
rect 1167 15 1173 21
rect 1263 39 1269 45
rect 1263 27 1269 33
rect 1263 15 1269 21
<< metal2 >>
rect -12 441 0 444
rect -12 435 -9 441
rect -3 435 0 441
rect -12 429 0 435
rect -12 423 -9 429
rect -3 423 0 429
rect -12 417 0 423
rect -12 411 -9 417
rect -3 411 0 417
rect -12 408 0 411
rect 12 441 24 444
rect 12 435 15 441
rect 21 435 24 441
rect 12 429 24 435
rect 12 423 15 429
rect 21 423 24 429
rect 12 417 24 423
rect 12 411 15 417
rect 21 411 24 417
rect -12 357 0 360
rect -12 351 -9 357
rect -3 351 0 357
rect -12 345 0 351
rect -12 339 -9 345
rect -3 339 0 345
rect -12 333 0 339
rect -12 327 -9 333
rect -3 327 0 333
rect -12 237 0 327
rect 12 357 24 411
rect 36 441 48 444
rect 36 435 39 441
rect 45 435 48 441
rect 36 429 48 435
rect 36 423 39 429
rect 45 423 48 429
rect 36 417 48 423
rect 36 411 39 417
rect 45 411 48 417
rect 36 408 48 411
rect 60 441 72 444
rect 60 435 63 441
rect 69 435 72 441
rect 60 429 72 435
rect 60 423 63 429
rect 69 423 72 429
rect 60 417 72 423
rect 60 411 63 417
rect 69 411 72 417
rect 36 393 48 396
rect 36 387 39 393
rect 45 387 48 393
rect 36 384 48 387
rect 12 351 15 357
rect 21 351 24 357
rect 12 345 24 351
rect 12 339 15 345
rect 21 339 24 345
rect 12 333 24 339
rect 12 327 15 333
rect 21 327 24 333
rect 12 324 24 327
rect 36 357 48 360
rect 36 351 39 357
rect 45 351 48 357
rect 36 345 48 351
rect 36 339 39 345
rect 45 339 48 345
rect 36 333 48 339
rect 36 327 39 333
rect 45 327 48 333
rect 12 309 24 312
rect 12 303 15 309
rect 21 303 24 309
rect 12 300 24 303
rect -12 231 -9 237
rect -3 231 0 237
rect -12 228 0 231
rect 12 228 24 240
rect 36 237 48 327
rect 60 357 72 411
rect 84 441 96 444
rect 84 435 87 441
rect 93 435 96 441
rect 84 429 96 435
rect 84 423 87 429
rect 93 423 96 429
rect 84 417 96 423
rect 84 411 87 417
rect 93 411 96 417
rect 84 408 96 411
rect 108 441 120 444
rect 108 435 111 441
rect 117 435 120 441
rect 108 429 120 435
rect 108 423 111 429
rect 117 423 120 429
rect 108 417 120 423
rect 108 411 111 417
rect 117 411 120 417
rect 84 393 96 396
rect 84 387 87 393
rect 93 387 96 393
rect 84 384 96 387
rect 60 351 63 357
rect 69 351 72 357
rect 60 345 72 351
rect 60 339 63 345
rect 69 339 72 345
rect 60 333 72 339
rect 60 327 63 333
rect 69 327 72 333
rect 60 324 72 327
rect 84 357 96 360
rect 84 351 87 357
rect 93 351 96 357
rect 84 345 96 351
rect 84 339 87 345
rect 93 339 96 345
rect 84 333 96 339
rect 84 327 87 333
rect 93 327 96 333
rect 60 309 72 312
rect 60 303 63 309
rect 69 303 72 309
rect 60 300 72 303
rect 36 231 39 237
rect 45 231 48 237
rect 36 228 48 231
rect 60 228 72 240
rect 84 237 96 327
rect 108 357 120 411
rect 132 441 144 444
rect 132 435 135 441
rect 141 435 144 441
rect 132 429 144 435
rect 132 423 135 429
rect 141 423 144 429
rect 132 417 144 423
rect 132 411 135 417
rect 141 411 144 417
rect 132 408 144 411
rect 156 441 168 444
rect 156 435 159 441
rect 165 435 168 441
rect 156 429 168 435
rect 156 423 159 429
rect 165 423 168 429
rect 156 417 168 423
rect 156 411 159 417
rect 165 411 168 417
rect 132 393 144 396
rect 132 387 135 393
rect 141 387 144 393
rect 132 384 144 387
rect 108 351 111 357
rect 117 351 120 357
rect 108 345 120 351
rect 108 339 111 345
rect 117 339 120 345
rect 108 333 120 339
rect 108 327 111 333
rect 117 327 120 333
rect 108 324 120 327
rect 132 357 144 360
rect 132 351 135 357
rect 141 351 144 357
rect 132 345 144 351
rect 132 339 135 345
rect 141 339 144 345
rect 132 333 144 339
rect 132 327 135 333
rect 141 327 144 333
rect 108 309 120 312
rect 108 303 111 309
rect 117 303 120 309
rect 108 300 120 303
rect 84 231 87 237
rect 93 231 96 237
rect 84 228 96 231
rect 132 237 144 327
rect 156 357 168 411
rect 180 441 192 444
rect 180 435 183 441
rect 189 435 192 441
rect 180 429 192 435
rect 180 423 183 429
rect 189 423 192 429
rect 180 417 192 423
rect 180 411 183 417
rect 189 411 192 417
rect 180 408 192 411
rect 204 441 216 444
rect 204 435 207 441
rect 213 435 216 441
rect 204 429 216 435
rect 204 423 207 429
rect 213 423 216 429
rect 204 417 216 423
rect 204 411 207 417
rect 213 411 216 417
rect 204 408 216 411
rect 252 441 264 444
rect 252 435 255 441
rect 261 435 264 441
rect 252 429 264 435
rect 252 423 255 429
rect 261 423 264 429
rect 252 417 264 423
rect 252 411 255 417
rect 261 411 264 417
rect 228 393 240 396
rect 228 387 231 393
rect 237 387 240 393
rect 228 384 240 387
rect 156 351 159 357
rect 165 351 168 357
rect 156 345 168 351
rect 156 339 159 345
rect 165 339 168 345
rect 156 333 168 339
rect 156 327 159 333
rect 165 327 168 333
rect 156 324 168 327
rect 180 357 192 360
rect 180 351 183 357
rect 189 351 192 357
rect 180 345 192 351
rect 180 339 183 345
rect 189 339 192 345
rect 180 333 192 339
rect 180 327 183 333
rect 189 327 192 333
rect 156 309 168 312
rect 156 303 159 309
rect 165 303 168 309
rect 156 300 168 303
rect 132 231 135 237
rect 141 231 144 237
rect 132 228 144 231
rect 180 237 192 327
rect 180 231 183 237
rect 189 231 192 237
rect 180 228 192 231
rect 204 357 216 360
rect 204 351 207 357
rect 213 351 216 357
rect 204 345 216 351
rect 204 339 207 345
rect 213 339 216 345
rect 204 333 216 339
rect 204 327 207 333
rect 213 327 216 333
rect -12 213 0 216
rect -12 207 -9 213
rect -3 207 0 213
rect -12 201 0 207
rect -12 195 -9 201
rect -3 195 0 201
rect -12 189 0 195
rect -12 183 -9 189
rect -3 183 0 189
rect -12 165 0 183
rect -12 159 -9 165
rect -3 159 0 165
rect -12 156 0 159
rect 36 213 48 216
rect 36 207 39 213
rect 45 207 48 213
rect 36 201 48 207
rect 36 195 39 201
rect 45 195 48 201
rect 36 189 48 195
rect 36 183 39 189
rect 45 183 48 189
rect 36 165 48 183
rect 36 159 39 165
rect 45 159 48 165
rect 36 156 48 159
rect 84 213 96 216
rect 84 207 87 213
rect 93 207 96 213
rect 84 201 96 207
rect 84 195 87 201
rect 93 195 96 201
rect 84 189 96 195
rect 84 183 87 189
rect 93 183 96 189
rect 84 165 96 183
rect 84 159 87 165
rect 93 159 96 165
rect 36 141 48 144
rect 36 135 39 141
rect 45 135 48 141
rect 12 69 24 72
rect 12 63 15 69
rect 21 63 24 69
rect 12 60 24 63
rect -12 45 0 48
rect -12 39 -9 45
rect -3 39 0 45
rect -12 33 0 39
rect -12 27 -9 33
rect -3 27 0 33
rect -12 21 0 27
rect -12 15 -9 21
rect -3 15 0 21
rect -12 12 0 15
rect 36 45 48 135
rect 60 69 72 72
rect 60 63 63 69
rect 69 63 72 69
rect 60 60 72 63
rect 36 39 39 45
rect 45 39 48 45
rect 36 33 48 39
rect 36 27 39 33
rect 45 27 48 33
rect 36 21 48 27
rect 36 15 39 21
rect 45 15 48 21
rect 36 12 48 15
rect 84 45 96 159
rect 132 213 144 216
rect 132 207 135 213
rect 141 207 144 213
rect 132 201 144 207
rect 132 195 135 201
rect 141 195 144 201
rect 132 189 144 195
rect 132 183 135 189
rect 141 183 144 189
rect 132 165 144 183
rect 132 159 135 165
rect 141 159 144 165
rect 132 156 144 159
rect 180 213 192 216
rect 180 207 183 213
rect 189 207 192 213
rect 180 201 192 207
rect 180 195 183 201
rect 189 195 192 201
rect 180 189 192 195
rect 180 183 183 189
rect 189 183 192 189
rect 180 165 192 183
rect 204 213 216 327
rect 252 357 264 411
rect 300 441 312 444
rect 300 435 303 441
rect 309 435 312 441
rect 300 429 312 435
rect 300 423 303 429
rect 309 423 312 429
rect 300 417 312 423
rect 300 411 303 417
rect 309 411 312 417
rect 300 408 312 411
rect 348 441 360 444
rect 348 435 351 441
rect 357 435 360 441
rect 348 429 360 435
rect 348 423 351 429
rect 357 423 360 429
rect 348 417 360 423
rect 348 411 351 417
rect 357 411 360 417
rect 276 393 288 396
rect 276 387 279 393
rect 285 387 288 393
rect 276 384 288 387
rect 324 393 336 396
rect 324 387 327 393
rect 333 387 336 393
rect 324 384 336 387
rect 252 351 255 357
rect 261 351 264 357
rect 252 345 264 351
rect 252 339 255 345
rect 261 339 264 345
rect 252 333 264 339
rect 252 327 255 333
rect 261 327 264 333
rect 252 324 264 327
rect 300 357 312 360
rect 300 351 303 357
rect 309 351 312 357
rect 300 345 312 351
rect 300 339 303 345
rect 309 339 312 345
rect 300 333 312 339
rect 300 327 303 333
rect 309 327 312 333
rect 300 324 312 327
rect 348 357 360 411
rect 396 441 408 444
rect 396 435 399 441
rect 405 435 408 441
rect 396 429 408 435
rect 396 423 399 429
rect 405 423 408 429
rect 396 417 408 423
rect 396 411 399 417
rect 405 411 408 417
rect 396 408 408 411
rect 420 441 432 444
rect 420 435 423 441
rect 429 435 432 441
rect 420 429 432 435
rect 420 423 423 429
rect 429 423 432 429
rect 420 417 432 423
rect 420 411 423 417
rect 429 411 432 417
rect 420 408 432 411
rect 468 441 480 444
rect 468 435 471 441
rect 477 435 480 441
rect 468 429 480 435
rect 468 423 471 429
rect 477 423 480 429
rect 468 417 480 423
rect 468 411 471 417
rect 477 411 480 417
rect 372 393 384 396
rect 372 387 375 393
rect 381 387 384 393
rect 372 384 384 387
rect 348 351 351 357
rect 357 351 360 357
rect 348 345 360 351
rect 348 339 351 345
rect 357 339 360 345
rect 348 333 360 339
rect 348 327 351 333
rect 357 327 360 333
rect 348 324 360 327
rect 396 357 408 360
rect 396 351 399 357
rect 405 351 408 357
rect 396 345 408 351
rect 396 339 399 345
rect 405 339 408 345
rect 396 333 408 339
rect 396 327 399 333
rect 405 327 408 333
rect 228 309 240 312
rect 228 303 231 309
rect 237 303 240 309
rect 228 300 240 303
rect 276 309 288 312
rect 276 303 279 309
rect 285 303 288 309
rect 276 300 288 303
rect 324 309 336 312
rect 324 303 327 309
rect 333 303 336 309
rect 324 300 336 303
rect 372 309 384 312
rect 372 303 375 309
rect 381 303 384 309
rect 372 300 384 303
rect 228 237 240 240
rect 228 231 231 237
rect 237 231 240 237
rect 228 228 240 231
rect 276 237 288 240
rect 276 231 279 237
rect 285 231 288 237
rect 276 228 288 231
rect 324 237 336 240
rect 324 231 327 237
rect 333 231 336 237
rect 324 228 336 231
rect 372 237 384 240
rect 372 231 375 237
rect 381 231 384 237
rect 372 228 384 231
rect 204 207 207 213
rect 213 207 216 213
rect 204 201 216 207
rect 204 195 207 201
rect 213 195 216 201
rect 204 189 216 195
rect 204 183 207 189
rect 213 183 216 189
rect 204 180 216 183
rect 300 213 312 216
rect 300 207 303 213
rect 309 207 312 213
rect 300 201 312 207
rect 300 195 303 201
rect 309 195 312 201
rect 300 189 312 195
rect 300 183 303 189
rect 309 183 312 189
rect 180 159 183 165
rect 189 159 192 165
rect 180 156 192 159
rect 132 141 144 144
rect 132 135 135 141
rect 141 135 144 141
rect 108 69 120 72
rect 108 63 111 69
rect 117 63 120 69
rect 108 60 120 63
rect 84 39 87 45
rect 93 39 96 45
rect 84 33 96 39
rect 84 27 87 33
rect 93 27 96 33
rect 84 21 96 27
rect 84 15 87 21
rect 93 15 96 21
rect 84 12 96 15
rect 132 45 144 135
rect 252 141 264 144
rect 252 135 255 141
rect 261 135 264 141
rect 156 69 168 72
rect 156 63 159 69
rect 165 63 168 69
rect 156 60 168 63
rect 228 69 240 72
rect 228 63 231 69
rect 237 63 240 69
rect 228 60 240 63
rect 132 39 135 45
rect 141 39 144 45
rect 132 33 144 39
rect 132 27 135 33
rect 141 27 144 33
rect 132 21 144 27
rect 132 15 135 21
rect 141 15 144 21
rect 132 12 144 15
rect 180 45 192 48
rect 180 39 183 45
rect 189 39 192 45
rect 180 33 192 39
rect 180 27 183 33
rect 189 27 192 33
rect 180 21 192 27
rect 180 15 183 21
rect 189 15 192 21
rect 180 12 192 15
rect 204 45 216 48
rect 204 39 207 45
rect 213 39 216 45
rect 204 33 216 39
rect 204 27 207 33
rect 213 27 216 33
rect 204 21 216 27
rect 204 15 207 21
rect 213 15 216 21
rect 204 12 216 15
rect 252 45 264 135
rect 300 117 312 183
rect 396 213 408 327
rect 396 207 399 213
rect 405 207 408 213
rect 396 201 408 207
rect 396 195 399 201
rect 405 195 408 201
rect 396 189 408 195
rect 396 183 399 189
rect 405 183 408 189
rect 396 180 408 183
rect 420 357 432 360
rect 420 351 423 357
rect 429 351 432 357
rect 420 345 432 351
rect 420 339 423 345
rect 429 339 432 345
rect 420 333 432 339
rect 420 327 423 333
rect 429 327 432 333
rect 420 237 432 327
rect 468 357 480 411
rect 516 441 528 444
rect 516 435 519 441
rect 525 435 528 441
rect 516 429 528 435
rect 516 423 519 429
rect 525 423 528 429
rect 516 417 528 423
rect 516 411 519 417
rect 525 411 528 417
rect 516 408 528 411
rect 564 441 576 444
rect 564 435 567 441
rect 573 435 576 441
rect 564 429 576 435
rect 564 423 567 429
rect 573 423 576 429
rect 564 417 576 423
rect 564 411 567 417
rect 573 411 576 417
rect 516 393 528 396
rect 516 387 519 393
rect 525 387 528 393
rect 516 384 528 387
rect 468 351 471 357
rect 477 351 480 357
rect 468 345 480 351
rect 468 339 471 345
rect 477 339 480 345
rect 468 333 480 339
rect 468 327 471 333
rect 477 327 480 333
rect 468 324 480 327
rect 516 357 528 360
rect 516 351 519 357
rect 525 351 528 357
rect 516 345 528 351
rect 516 339 519 345
rect 525 339 528 345
rect 516 333 528 339
rect 516 327 519 333
rect 525 327 528 333
rect 516 324 528 327
rect 564 357 576 411
rect 612 441 624 444
rect 612 435 615 441
rect 621 435 624 441
rect 612 429 624 435
rect 612 423 615 429
rect 621 423 624 429
rect 612 417 624 423
rect 612 411 615 417
rect 621 411 624 417
rect 612 408 624 411
rect 636 441 648 444
rect 636 435 639 441
rect 645 435 648 441
rect 636 429 648 435
rect 636 423 639 429
rect 645 423 648 429
rect 636 417 648 423
rect 636 411 639 417
rect 645 411 648 417
rect 636 408 648 411
rect 828 441 840 444
rect 828 435 831 441
rect 837 435 840 441
rect 828 429 840 435
rect 828 423 831 429
rect 837 423 840 429
rect 828 417 840 423
rect 828 411 831 417
rect 837 411 840 417
rect 636 393 648 396
rect 636 387 639 393
rect 645 387 648 393
rect 564 351 567 357
rect 573 351 576 357
rect 564 345 576 351
rect 564 339 567 345
rect 573 339 576 345
rect 564 333 576 339
rect 564 327 567 333
rect 573 327 576 333
rect 564 324 576 327
rect 612 357 624 360
rect 612 351 615 357
rect 621 351 624 357
rect 612 345 624 351
rect 612 339 615 345
rect 621 339 624 345
rect 612 333 624 339
rect 612 327 615 333
rect 621 327 624 333
rect 444 309 456 312
rect 444 303 447 309
rect 453 303 456 309
rect 444 300 456 303
rect 492 309 504 312
rect 492 303 495 309
rect 501 303 504 309
rect 492 300 504 303
rect 540 309 552 312
rect 540 303 543 309
rect 549 303 552 309
rect 540 300 552 303
rect 588 309 600 312
rect 588 303 591 309
rect 597 303 600 309
rect 588 300 600 303
rect 420 231 423 237
rect 429 231 432 237
rect 420 213 432 231
rect 444 237 456 240
rect 444 231 447 237
rect 453 231 456 237
rect 444 228 456 231
rect 492 237 504 240
rect 492 231 495 237
rect 501 231 504 237
rect 492 228 504 231
rect 540 237 552 240
rect 540 231 543 237
rect 549 231 552 237
rect 540 228 552 231
rect 588 237 600 240
rect 588 231 591 237
rect 597 231 600 237
rect 588 228 600 231
rect 420 207 423 213
rect 429 207 432 213
rect 420 201 432 207
rect 420 195 423 201
rect 429 195 432 201
rect 420 189 432 195
rect 420 183 423 189
rect 429 183 432 189
rect 420 180 432 183
rect 516 213 528 216
rect 516 207 519 213
rect 525 207 528 213
rect 516 201 528 207
rect 516 195 519 201
rect 525 195 528 201
rect 516 189 528 195
rect 516 183 519 189
rect 525 183 528 189
rect 300 111 303 117
rect 309 111 312 117
rect 276 69 288 72
rect 276 63 279 69
rect 285 63 288 69
rect 276 60 288 63
rect 252 39 255 45
rect 261 39 264 45
rect 252 33 264 39
rect 252 27 255 33
rect 261 27 264 33
rect 252 21 264 27
rect 252 15 255 21
rect 261 15 264 21
rect 252 12 264 15
rect 300 45 312 111
rect 348 141 360 144
rect 348 135 351 141
rect 357 135 360 141
rect 324 69 336 72
rect 324 63 327 69
rect 333 63 336 69
rect 324 60 336 63
rect 300 39 303 45
rect 309 39 312 45
rect 300 33 312 39
rect 300 27 303 33
rect 309 27 312 33
rect 300 21 312 27
rect 300 15 303 21
rect 309 15 312 21
rect 300 12 312 15
rect 348 45 360 135
rect 516 93 528 183
rect 612 213 624 327
rect 612 207 615 213
rect 621 207 624 213
rect 612 201 624 207
rect 612 195 615 201
rect 621 195 624 201
rect 612 189 624 195
rect 612 183 615 189
rect 621 183 624 189
rect 612 180 624 183
rect 636 357 648 387
rect 636 351 639 357
rect 645 351 648 357
rect 636 345 648 351
rect 636 339 639 345
rect 645 339 648 345
rect 636 333 648 339
rect 636 327 639 333
rect 645 327 648 333
rect 636 309 648 327
rect 828 357 840 411
rect 828 351 831 357
rect 837 351 840 357
rect 828 345 840 351
rect 828 339 831 345
rect 837 339 840 345
rect 828 333 840 339
rect 828 327 831 333
rect 837 327 840 333
rect 828 324 840 327
rect 852 441 864 444
rect 852 435 855 441
rect 861 435 864 441
rect 852 429 864 435
rect 852 423 855 429
rect 861 423 864 429
rect 852 417 864 423
rect 852 411 855 417
rect 861 411 864 417
rect 852 357 864 411
rect 1044 441 1056 444
rect 1044 435 1047 441
rect 1053 435 1056 441
rect 1044 429 1056 435
rect 1044 423 1047 429
rect 1053 423 1056 429
rect 1044 417 1056 423
rect 1044 411 1047 417
rect 1053 411 1056 417
rect 852 351 855 357
rect 861 351 864 357
rect 852 345 864 351
rect 852 339 855 345
rect 861 339 864 345
rect 852 333 864 339
rect 852 327 855 333
rect 861 327 864 333
rect 852 324 864 327
rect 900 393 912 396
rect 900 387 903 393
rect 909 387 912 393
rect 636 303 639 309
rect 645 303 648 309
rect 636 213 648 303
rect 660 309 672 312
rect 660 303 663 309
rect 669 303 672 309
rect 660 300 672 303
rect 708 309 720 312
rect 708 303 711 309
rect 717 303 720 309
rect 708 300 720 303
rect 756 309 768 312
rect 756 303 759 309
rect 765 303 768 309
rect 756 300 768 303
rect 804 309 816 312
rect 804 303 807 309
rect 813 303 816 309
rect 804 300 816 303
rect 828 309 840 312
rect 828 303 831 309
rect 837 303 840 309
rect 660 237 672 240
rect 660 231 663 237
rect 669 231 672 237
rect 660 228 672 231
rect 708 237 720 240
rect 708 231 711 237
rect 717 231 720 237
rect 708 228 720 231
rect 756 237 768 240
rect 756 231 759 237
rect 765 231 768 237
rect 756 228 768 231
rect 804 237 816 240
rect 804 231 807 237
rect 813 231 816 237
rect 804 228 816 231
rect 636 207 639 213
rect 645 207 648 213
rect 636 201 648 207
rect 636 195 639 201
rect 645 195 648 201
rect 636 189 648 195
rect 636 183 639 189
rect 645 183 648 189
rect 636 180 648 183
rect 732 213 744 216
rect 732 207 735 213
rect 741 207 744 213
rect 732 201 744 207
rect 732 195 735 201
rect 741 195 744 201
rect 732 189 744 195
rect 732 183 735 189
rect 741 183 744 189
rect 516 87 519 93
rect 525 87 528 93
rect 372 69 384 72
rect 372 63 375 69
rect 381 63 384 69
rect 372 60 384 63
rect 444 69 456 72
rect 444 63 447 69
rect 453 63 456 69
rect 444 60 456 63
rect 492 69 504 72
rect 492 63 495 69
rect 501 63 504 69
rect 492 60 504 63
rect 348 39 351 45
rect 357 39 360 45
rect 348 33 360 39
rect 348 27 351 33
rect 357 27 360 33
rect 348 21 360 27
rect 348 15 351 21
rect 357 15 360 21
rect 348 12 360 15
rect 396 45 408 48
rect 396 39 399 45
rect 405 39 408 45
rect 396 33 408 39
rect 396 27 399 33
rect 405 27 408 33
rect 396 21 408 27
rect 396 15 399 21
rect 405 15 408 21
rect 396 12 408 15
rect 420 45 432 48
rect 420 39 423 45
rect 429 39 432 45
rect 420 33 432 39
rect 420 27 423 33
rect 429 27 432 33
rect 420 21 432 27
rect 420 15 423 21
rect 429 15 432 21
rect 420 12 432 15
rect 516 45 528 87
rect 540 69 552 72
rect 540 63 543 69
rect 549 63 552 69
rect 540 60 552 63
rect 588 69 600 72
rect 588 63 591 69
rect 597 63 600 69
rect 588 60 600 63
rect 660 69 672 72
rect 660 63 663 69
rect 669 63 672 69
rect 660 60 672 63
rect 708 69 720 72
rect 708 63 711 69
rect 717 63 720 69
rect 708 60 720 63
rect 516 39 519 45
rect 525 39 528 45
rect 516 33 528 39
rect 516 27 519 33
rect 525 27 528 33
rect 516 21 528 27
rect 516 15 519 21
rect 525 15 528 21
rect 516 12 528 15
rect 612 45 624 48
rect 612 39 615 45
rect 621 39 624 45
rect 612 33 624 39
rect 612 27 615 33
rect 621 27 624 33
rect 612 21 624 27
rect 612 15 615 21
rect 621 15 624 21
rect 612 12 624 15
rect 636 45 648 48
rect 636 39 639 45
rect 645 39 648 45
rect 636 33 648 39
rect 636 27 639 33
rect 645 27 648 33
rect 636 21 648 27
rect 636 15 639 21
rect 645 15 648 21
rect 636 12 648 15
rect 732 45 744 183
rect 828 213 840 303
rect 900 309 912 387
rect 1044 357 1056 411
rect 1044 351 1047 357
rect 1053 351 1056 357
rect 1044 345 1056 351
rect 1044 339 1047 345
rect 1053 339 1056 345
rect 1044 333 1056 339
rect 1044 327 1047 333
rect 1053 327 1056 333
rect 1044 324 1056 327
rect 900 303 903 309
rect 909 303 912 309
rect 900 240 912 303
rect 864 237 912 240
rect 864 231 867 237
rect 873 231 912 237
rect 864 228 912 231
rect 924 237 936 240
rect 924 231 927 237
rect 933 231 936 237
rect 924 228 936 231
rect 972 237 984 240
rect 972 231 975 237
rect 981 231 984 237
rect 972 228 984 231
rect 1020 237 1032 240
rect 1020 231 1023 237
rect 1029 231 1032 237
rect 1020 228 1032 231
rect 1092 237 1104 240
rect 1092 231 1095 237
rect 1101 231 1104 237
rect 1092 228 1104 231
rect 1140 237 1152 240
rect 1140 231 1143 237
rect 1149 231 1152 237
rect 1140 228 1152 231
rect 1188 237 1200 240
rect 1188 231 1191 237
rect 1197 231 1200 237
rect 1188 228 1200 231
rect 1236 237 1248 240
rect 1236 231 1239 237
rect 1245 231 1248 237
rect 1236 228 1248 231
rect 828 207 831 213
rect 837 207 840 213
rect 828 201 840 207
rect 828 195 831 201
rect 837 195 840 201
rect 828 189 840 195
rect 828 183 831 189
rect 837 183 840 189
rect 828 180 840 183
rect 852 213 864 216
rect 852 207 855 213
rect 861 207 864 213
rect 852 201 864 207
rect 852 195 855 201
rect 861 195 864 201
rect 852 189 864 195
rect 852 183 855 189
rect 861 183 864 189
rect 852 180 864 183
rect 876 213 888 216
rect 876 207 879 213
rect 885 207 888 213
rect 876 201 888 207
rect 876 195 879 201
rect 885 195 888 201
rect 876 189 888 195
rect 876 183 879 189
rect 885 183 888 189
rect 876 180 888 183
rect 900 213 912 228
rect 900 207 903 213
rect 909 207 912 213
rect 900 201 912 207
rect 900 195 903 201
rect 909 195 912 201
rect 900 189 912 195
rect 900 183 903 189
rect 909 183 912 189
rect 900 180 912 183
rect 1044 213 1056 216
rect 1044 207 1047 213
rect 1053 207 1056 213
rect 1044 201 1056 207
rect 1044 195 1047 201
rect 1053 195 1056 201
rect 1044 189 1056 195
rect 1044 183 1047 189
rect 1053 183 1056 189
rect 756 69 768 72
rect 756 63 759 69
rect 765 63 768 69
rect 756 60 768 63
rect 804 69 816 72
rect 804 63 807 69
rect 813 63 816 69
rect 804 60 816 63
rect 876 69 888 72
rect 876 63 879 69
rect 885 63 888 69
rect 876 60 888 63
rect 924 69 936 72
rect 924 63 927 69
rect 933 63 936 69
rect 924 60 936 63
rect 972 69 984 72
rect 972 63 975 69
rect 981 63 984 69
rect 972 60 984 63
rect 1020 69 1032 72
rect 1020 63 1023 69
rect 1029 63 1032 69
rect 1020 60 1032 63
rect 732 39 735 45
rect 741 39 744 45
rect 732 33 744 39
rect 732 27 735 33
rect 741 27 744 33
rect 732 21 744 27
rect 732 15 735 21
rect 741 15 744 21
rect 732 12 744 15
rect 828 45 840 48
rect 828 39 831 45
rect 837 39 840 45
rect 828 33 840 39
rect 828 27 831 33
rect 837 27 840 33
rect 828 21 840 27
rect 828 15 831 21
rect 837 15 840 21
rect 828 12 840 15
rect 852 45 864 48
rect 852 39 855 45
rect 861 39 864 45
rect 852 33 864 39
rect 852 27 855 33
rect 861 27 864 33
rect 852 21 864 27
rect 852 15 855 21
rect 861 15 864 21
rect 852 12 864 15
rect 1044 45 1056 183
rect 1068 213 1080 216
rect 1068 207 1071 213
rect 1077 207 1080 213
rect 1068 201 1080 207
rect 1068 195 1071 201
rect 1077 195 1080 201
rect 1068 189 1080 195
rect 1068 183 1071 189
rect 1077 183 1080 189
rect 1068 180 1080 183
rect 1164 213 1176 216
rect 1164 207 1167 213
rect 1173 207 1176 213
rect 1164 201 1176 207
rect 1164 195 1167 201
rect 1173 195 1176 201
rect 1164 189 1176 195
rect 1164 183 1167 189
rect 1173 183 1176 189
rect 1092 69 1104 72
rect 1092 63 1095 69
rect 1101 63 1104 69
rect 1092 60 1104 63
rect 1140 69 1152 72
rect 1140 63 1143 69
rect 1149 63 1152 69
rect 1140 60 1152 63
rect 1044 39 1047 45
rect 1053 39 1056 45
rect 1044 33 1056 39
rect 1044 27 1047 33
rect 1053 27 1056 33
rect 1044 21 1056 27
rect 1044 15 1047 21
rect 1053 15 1056 21
rect 1044 12 1056 15
rect 1068 45 1080 48
rect 1068 39 1071 45
rect 1077 39 1080 45
rect 1068 33 1080 39
rect 1068 27 1071 33
rect 1077 27 1080 33
rect 1068 21 1080 27
rect 1068 15 1071 21
rect 1077 15 1080 21
rect 1068 12 1080 15
rect 1164 45 1176 183
rect 1260 213 1272 216
rect 1260 207 1263 213
rect 1269 207 1272 213
rect 1260 201 1272 207
rect 1260 195 1263 201
rect 1269 195 1272 201
rect 1260 189 1272 195
rect 1260 183 1263 189
rect 1269 183 1272 189
rect 1260 180 1272 183
rect 1188 69 1200 72
rect 1188 63 1191 69
rect 1197 63 1200 69
rect 1188 60 1200 63
rect 1236 69 1248 72
rect 1236 63 1239 69
rect 1245 63 1248 69
rect 1236 60 1248 63
rect 1164 39 1167 45
rect 1173 39 1176 45
rect 1164 33 1176 39
rect 1164 27 1167 33
rect 1173 27 1176 33
rect 1164 21 1176 27
rect 1164 15 1167 21
rect 1173 15 1176 21
rect 1164 12 1176 15
rect 1260 45 1272 48
rect 1260 39 1263 45
rect 1269 39 1272 45
rect 1260 33 1272 39
rect 1260 27 1263 33
rect 1269 27 1272 33
rect 1260 21 1272 27
rect 1260 15 1263 21
rect 1269 15 1272 21
rect 1260 12 1272 15
<< via2 >>
rect -9 435 -3 441
rect -9 423 -3 429
rect -9 411 -3 417
rect -9 327 -3 333
rect 39 435 45 441
rect 39 423 45 429
rect 39 411 45 417
rect 39 387 45 393
rect 15 351 21 357
rect 39 327 45 333
rect 15 303 21 309
rect 87 435 93 441
rect 87 423 93 429
rect 87 411 93 417
rect 87 387 93 393
rect 63 351 69 357
rect 87 327 93 333
rect 63 303 69 309
rect 135 435 141 441
rect 135 423 141 429
rect 135 411 141 417
rect 135 387 141 393
rect 111 351 117 357
rect 135 327 141 333
rect 111 303 117 309
rect 183 435 189 441
rect 183 423 189 429
rect 183 411 189 417
rect 207 435 213 441
rect 207 423 213 429
rect 207 411 213 417
rect 231 387 237 393
rect 159 351 165 357
rect 183 327 189 333
rect 159 303 165 309
rect 207 327 213 333
rect -9 159 -3 165
rect 39 159 45 165
rect 87 159 93 165
rect 39 135 45 141
rect 15 63 21 69
rect -9 39 -3 45
rect -9 27 -3 33
rect -9 15 -3 21
rect 63 63 69 69
rect 135 159 141 165
rect 303 435 309 441
rect 303 423 309 429
rect 303 411 309 417
rect 279 387 285 393
rect 327 387 333 393
rect 255 351 261 357
rect 303 327 309 333
rect 399 435 405 441
rect 399 423 405 429
rect 399 411 405 417
rect 423 435 429 441
rect 423 423 429 429
rect 423 411 429 417
rect 375 387 381 393
rect 351 351 357 357
rect 399 327 405 333
rect 231 303 237 309
rect 279 303 285 309
rect 327 303 333 309
rect 375 303 381 309
rect 231 231 237 237
rect 279 231 285 237
rect 327 231 333 237
rect 375 231 381 237
rect 183 159 189 165
rect 135 135 141 141
rect 111 63 117 69
rect 255 135 261 141
rect 159 63 165 69
rect 231 63 237 69
rect 183 39 189 45
rect 183 27 189 33
rect 183 15 189 21
rect 207 39 213 45
rect 207 27 213 33
rect 207 15 213 21
rect 423 327 429 333
rect 519 435 525 441
rect 519 423 525 429
rect 519 411 525 417
rect 519 387 525 393
rect 471 351 477 357
rect 519 327 525 333
rect 615 435 621 441
rect 615 423 621 429
rect 615 411 621 417
rect 639 435 645 441
rect 639 423 645 429
rect 639 411 645 417
rect 567 351 573 357
rect 615 327 621 333
rect 447 303 453 309
rect 495 303 501 309
rect 543 303 549 309
rect 591 303 597 309
rect 423 231 429 237
rect 447 231 453 237
rect 495 231 501 237
rect 543 231 549 237
rect 591 231 597 237
rect 303 111 309 117
rect 279 63 285 69
rect 351 135 357 141
rect 327 63 333 69
rect 639 303 645 309
rect 663 303 669 309
rect 711 303 717 309
rect 759 303 765 309
rect 807 303 813 309
rect 663 231 669 237
rect 711 231 717 237
rect 759 231 765 237
rect 807 231 813 237
rect 519 87 525 93
rect 375 63 381 69
rect 447 63 453 69
rect 495 63 501 69
rect 399 39 405 45
rect 399 27 405 33
rect 399 15 405 21
rect 423 39 429 45
rect 423 27 429 33
rect 423 15 429 21
rect 543 63 549 69
rect 591 63 597 69
rect 663 63 669 69
rect 711 63 717 69
rect 615 39 621 45
rect 615 27 621 33
rect 615 15 621 21
rect 639 39 645 45
rect 639 27 645 33
rect 639 15 645 21
rect 927 231 933 237
rect 975 231 981 237
rect 1023 231 1029 237
rect 1095 231 1101 237
rect 1143 231 1149 237
rect 1191 231 1197 237
rect 1239 231 1245 237
rect 759 63 765 69
rect 807 63 813 69
rect 879 63 885 69
rect 927 63 933 69
rect 975 63 981 69
rect 1023 63 1029 69
rect 831 39 837 45
rect 831 27 837 33
rect 831 15 837 21
rect 855 39 861 45
rect 855 27 861 33
rect 855 15 861 21
rect 1071 207 1077 213
rect 1095 63 1101 69
rect 1143 63 1149 69
rect 1071 39 1077 45
rect 1071 27 1077 33
rect 1071 15 1077 21
rect 1263 207 1269 213
rect 1191 63 1197 69
rect 1239 63 1245 69
rect 1263 39 1269 45
rect 1263 27 1269 33
rect 1263 15 1269 21
<< metal3 >>
rect -24 441 1068 444
rect -24 435 -9 441
rect -3 435 39 441
rect 45 435 87 441
rect 93 435 135 441
rect 141 435 183 441
rect 189 435 207 441
rect 213 435 303 441
rect 309 435 399 441
rect 405 435 423 441
rect 429 435 519 441
rect 525 435 615 441
rect 621 435 639 441
rect 645 435 1068 441
rect -24 429 1068 435
rect -24 423 -9 429
rect -3 423 39 429
rect 45 423 87 429
rect 93 423 135 429
rect 141 423 183 429
rect 189 423 207 429
rect 213 423 303 429
rect 309 423 399 429
rect 405 423 423 429
rect 429 423 519 429
rect 525 423 615 429
rect 621 423 639 429
rect 645 423 1068 429
rect -24 417 1068 423
rect -24 411 -9 417
rect -3 411 39 417
rect 45 411 87 417
rect 93 411 135 417
rect 141 411 183 417
rect 189 411 207 417
rect 213 411 303 417
rect 309 411 399 417
rect 405 411 423 417
rect 429 411 519 417
rect 525 411 615 417
rect 621 411 639 417
rect 645 411 1068 417
rect -24 408 1068 411
rect -24 393 1068 396
rect -24 387 39 393
rect 45 387 87 393
rect 93 387 135 393
rect 141 387 231 393
rect 237 387 279 393
rect 285 387 303 393
rect 309 387 327 393
rect 333 387 375 393
rect 381 387 519 393
rect 525 387 1068 393
rect -24 384 1068 387
rect 12 357 168 360
rect 12 351 15 357
rect 21 351 63 357
rect 69 351 111 357
rect 117 351 159 357
rect 165 351 168 357
rect 12 348 168 351
rect 252 357 360 360
rect 252 351 255 357
rect 261 351 351 357
rect 357 351 360 357
rect 252 348 360 351
rect 468 357 576 360
rect 468 351 471 357
rect 477 351 567 357
rect 573 351 576 357
rect 468 348 576 351
rect -12 333 192 336
rect -12 327 -9 333
rect -3 327 39 333
rect 45 327 87 333
rect 93 327 135 333
rect 141 327 183 333
rect 189 327 192 333
rect -12 324 192 327
rect 204 333 408 336
rect 204 327 207 333
rect 213 327 303 333
rect 309 327 399 333
rect 405 327 408 333
rect 204 324 408 327
rect 420 333 624 336
rect 420 327 423 333
rect 429 327 519 333
rect 525 327 615 333
rect 621 327 624 333
rect 420 324 624 327
rect -24 309 1068 312
rect -24 303 15 309
rect 21 303 63 309
rect 69 303 111 309
rect 117 303 159 309
rect 165 303 231 309
rect 237 303 279 309
rect 285 303 327 309
rect 333 303 375 309
rect 381 303 447 309
rect 453 303 495 309
rect 501 303 543 309
rect 549 303 591 309
rect 597 303 639 309
rect 645 303 663 309
rect 669 303 711 309
rect 717 303 759 309
rect 765 303 807 309
rect 813 303 855 309
rect 861 303 1068 309
rect -24 300 1068 303
rect 216 237 1284 240
rect 216 231 231 237
rect 237 231 279 237
rect 285 231 327 237
rect 333 231 375 237
rect 381 231 423 237
rect 429 231 447 237
rect 453 231 495 237
rect 501 231 543 237
rect 549 231 591 237
rect 597 231 663 237
rect 669 231 711 237
rect 717 231 759 237
rect 765 231 807 237
rect 813 231 927 237
rect 933 231 975 237
rect 981 231 1023 237
rect 1029 231 1095 237
rect 1101 231 1143 237
rect 1149 231 1191 237
rect 1197 231 1239 237
rect 1245 231 1284 237
rect 216 228 1284 231
rect 852 213 864 216
rect 852 207 855 213
rect 861 207 864 213
rect 852 201 864 207
rect 852 195 855 201
rect 861 195 864 201
rect 852 189 864 195
rect 852 183 855 189
rect 861 183 864 189
rect 852 180 864 183
rect 876 213 888 216
rect 876 207 879 213
rect 885 207 888 213
rect 876 201 888 207
rect 1068 213 1284 216
rect 1068 207 1071 213
rect 1077 207 1263 213
rect 1269 207 1284 213
rect 1068 204 1284 207
rect 876 195 879 201
rect 885 195 888 201
rect 876 189 888 195
rect 876 183 879 189
rect 885 183 888 189
rect 876 180 888 183
rect -24 165 1284 168
rect -24 159 -9 165
rect -3 159 15 165
rect 21 159 39 165
rect 45 159 63 165
rect 69 159 87 165
rect 93 159 111 165
rect 117 159 135 165
rect 141 159 159 165
rect 165 159 183 165
rect 189 159 231 165
rect 237 159 375 165
rect 381 159 1284 165
rect -24 156 1284 159
rect -24 141 1284 144
rect -24 135 39 141
rect 45 135 135 141
rect 141 135 255 141
rect 261 135 351 141
rect 357 135 1284 141
rect -24 132 1284 135
rect -24 117 1284 120
rect -24 111 303 117
rect 309 111 1284 117
rect -24 108 1284 111
rect -24 93 1284 96
rect -24 87 279 93
rect 285 87 327 93
rect 333 87 447 93
rect 453 87 495 93
rect 501 87 519 93
rect 525 87 543 93
rect 549 87 591 93
rect 597 87 663 93
rect 669 87 711 93
rect 717 87 759 93
rect 765 87 807 93
rect 813 87 879 93
rect 885 87 927 93
rect 933 87 975 93
rect 981 87 1023 93
rect 1029 87 1095 93
rect 1101 87 1143 93
rect 1149 87 1191 93
rect 1197 87 1239 93
rect 1245 87 1284 93
rect -24 84 1284 87
rect 12 69 24 72
rect 12 63 15 69
rect 21 63 24 69
rect 12 60 24 63
rect 60 69 72 72
rect 60 63 63 69
rect 69 63 72 69
rect 60 60 72 63
rect 108 69 120 72
rect 108 63 111 69
rect 117 63 120 69
rect 108 60 120 63
rect 156 69 168 72
rect 156 63 159 69
rect 165 63 168 69
rect 156 60 168 63
rect 228 69 240 72
rect 228 63 231 69
rect 237 63 240 69
rect 228 60 240 63
rect 276 69 288 72
rect 276 63 279 69
rect 285 63 288 69
rect 276 60 288 63
rect 324 69 336 72
rect 324 63 327 69
rect 333 63 336 69
rect 324 60 336 63
rect 372 69 384 72
rect 372 63 375 69
rect 381 63 384 69
rect 372 60 384 63
rect 444 69 456 72
rect 444 63 447 69
rect 453 63 456 69
rect 444 60 456 63
rect 492 69 504 72
rect 492 63 495 69
rect 501 63 504 69
rect 492 60 504 63
rect 540 69 552 72
rect 540 63 543 69
rect 549 63 552 69
rect 540 60 552 63
rect 588 69 600 72
rect 588 63 591 69
rect 597 63 600 69
rect 588 60 600 63
rect 660 69 672 72
rect 660 63 663 69
rect 669 63 672 69
rect 660 60 672 63
rect 708 69 720 72
rect 708 63 711 69
rect 717 63 720 69
rect 708 60 720 63
rect 756 69 768 72
rect 756 63 759 69
rect 765 63 768 69
rect 756 60 768 63
rect 804 69 816 72
rect 804 63 807 69
rect 813 63 816 69
rect 804 60 816 63
rect 876 69 888 72
rect 876 63 879 69
rect 885 63 888 69
rect 876 60 888 63
rect 924 69 936 72
rect 924 63 927 69
rect 933 63 936 69
rect 924 60 936 63
rect 972 69 984 72
rect 972 63 975 69
rect 981 63 984 69
rect 972 60 984 63
rect 1020 69 1032 72
rect 1020 63 1023 69
rect 1029 63 1032 69
rect 1020 60 1032 63
rect 1092 69 1104 72
rect 1092 63 1095 69
rect 1101 63 1104 69
rect 1092 60 1104 63
rect 1140 69 1152 72
rect 1140 63 1143 69
rect 1149 63 1152 69
rect 1140 60 1152 63
rect 1188 69 1200 72
rect 1188 63 1191 69
rect 1197 63 1200 69
rect 1188 60 1200 63
rect 1236 69 1248 72
rect 1236 63 1239 69
rect 1245 63 1248 69
rect 1236 60 1248 63
rect -24 45 1284 48
rect -24 39 -9 45
rect -3 39 183 45
rect 189 39 207 45
rect 213 39 399 45
rect 405 39 423 45
rect 429 39 615 45
rect 621 39 639 45
rect 645 39 831 45
rect 837 39 855 45
rect 861 39 1071 45
rect 1077 39 1263 45
rect 1269 39 1284 45
rect -24 33 1284 39
rect -24 27 -9 33
rect -3 27 183 33
rect 189 27 207 33
rect 213 27 399 33
rect 405 27 423 33
rect 429 27 615 33
rect 621 27 639 33
rect 645 27 831 33
rect 837 27 855 33
rect 861 27 1071 33
rect 1077 27 1263 33
rect 1269 27 1284 33
rect -24 21 1284 27
rect -24 15 -9 21
rect -3 15 183 21
rect 189 15 207 21
rect 213 15 399 21
rect 405 15 423 21
rect 429 15 615 21
rect 621 15 639 21
rect 645 15 831 21
rect 837 15 855 21
rect 861 15 1071 21
rect 1077 15 1263 21
rect 1269 15 1284 21
rect -24 12 1284 15
<< via3 >>
rect 303 387 309 393
rect 303 327 309 333
rect 855 303 861 309
rect 855 207 861 213
rect 855 195 861 201
rect 855 183 861 189
rect 879 207 885 213
rect 879 195 885 201
rect 879 183 885 189
rect 15 159 21 165
rect 63 159 69 165
rect 111 159 117 165
rect 159 159 165 165
rect 231 159 237 165
rect 375 159 381 165
rect 279 87 285 93
rect 327 87 333 93
rect 447 87 453 93
rect 495 87 501 93
rect 543 87 549 93
rect 591 87 597 93
rect 663 87 669 93
rect 711 87 717 93
rect 759 87 765 93
rect 807 87 813 93
rect 879 87 885 93
rect 927 87 933 93
rect 975 87 981 93
rect 1023 87 1029 93
rect 1095 87 1101 93
rect 1143 87 1149 93
rect 1191 87 1197 93
rect 1239 87 1245 93
rect 15 63 21 69
rect 63 63 69 69
rect 111 63 117 69
rect 159 63 165 69
rect 231 63 237 69
rect 279 63 285 69
rect 327 63 333 69
rect 375 63 381 69
rect 447 63 453 69
rect 495 63 501 69
rect 543 63 549 69
rect 591 63 597 69
rect 663 63 669 69
rect 711 63 717 69
rect 759 63 765 69
rect 807 63 813 69
rect 879 63 885 69
rect 927 63 933 69
rect 975 63 981 69
rect 1023 63 1029 69
rect 1095 63 1101 69
rect 1143 63 1149 69
rect 1191 63 1197 69
rect 1239 63 1245 69
<< metal4 >>
rect 852 420 864 444
rect 300 393 312 396
rect 300 387 303 393
rect 309 387 312 393
rect 300 333 312 387
rect 300 327 303 333
rect 309 327 312 333
rect 300 324 312 327
rect 852 309 864 312
rect 852 303 855 309
rect 861 303 864 309
rect 192 252 204 288
rect 408 252 420 288
rect 624 252 636 288
rect 852 213 864 303
rect 852 207 855 213
rect 861 207 864 213
rect 852 201 864 207
rect 852 195 855 201
rect 861 195 864 201
rect 852 189 864 195
rect 852 183 855 189
rect 861 183 864 189
rect 852 180 864 183
rect 876 213 888 216
rect 876 207 879 213
rect 885 207 888 213
rect 876 201 888 207
rect 876 195 879 201
rect 885 195 888 201
rect 876 189 888 195
rect 876 183 879 189
rect 885 183 888 189
rect 12 165 24 168
rect 12 159 15 165
rect 21 159 24 165
rect 12 69 24 159
rect 12 63 15 69
rect 21 63 24 69
rect 12 60 24 63
rect 60 165 72 168
rect 60 159 63 165
rect 69 159 72 165
rect 60 69 72 159
rect 60 63 63 69
rect 69 63 72 69
rect 60 60 72 63
rect 108 165 120 168
rect 108 159 111 165
rect 117 159 120 165
rect 108 69 120 159
rect 108 63 111 69
rect 117 63 120 69
rect 108 60 120 63
rect 156 165 168 168
rect 156 159 159 165
rect 165 159 168 165
rect 156 69 168 159
rect 156 63 159 69
rect 165 63 168 69
rect 156 60 168 63
rect 228 165 240 168
rect 228 159 231 165
rect 237 159 240 165
rect 228 69 240 159
rect 372 165 384 168
rect 372 159 375 165
rect 381 159 384 165
rect 228 63 231 69
rect 237 63 240 69
rect 228 60 240 63
rect 276 93 288 96
rect 276 87 279 93
rect 285 87 288 93
rect 276 69 288 87
rect 276 63 279 69
rect 285 63 288 69
rect 276 60 288 63
rect 324 93 336 96
rect 324 87 327 93
rect 333 87 336 93
rect 324 69 336 87
rect 324 63 327 69
rect 333 63 336 69
rect 324 60 336 63
rect 372 69 384 159
rect 372 63 375 69
rect 381 63 384 69
rect 372 60 384 63
rect 444 93 456 96
rect 444 87 447 93
rect 453 87 456 93
rect 444 69 456 87
rect 444 63 447 69
rect 453 63 456 69
rect 444 60 456 63
rect 492 93 504 96
rect 492 87 495 93
rect 501 87 504 93
rect 492 69 504 87
rect 492 63 495 69
rect 501 63 504 69
rect 492 60 504 63
rect 540 93 552 96
rect 540 87 543 93
rect 549 87 552 93
rect 540 69 552 87
rect 540 63 543 69
rect 549 63 552 69
rect 540 60 552 63
rect 588 93 600 96
rect 588 87 591 93
rect 597 87 600 93
rect 588 69 600 87
rect 588 63 591 69
rect 597 63 600 69
rect 588 60 600 63
rect 660 93 672 96
rect 660 87 663 93
rect 669 87 672 93
rect 660 69 672 87
rect 660 63 663 69
rect 669 63 672 69
rect 660 60 672 63
rect 708 93 720 96
rect 708 87 711 93
rect 717 87 720 93
rect 708 69 720 87
rect 708 63 711 69
rect 717 63 720 69
rect 708 60 720 63
rect 756 93 768 96
rect 756 87 759 93
rect 765 87 768 93
rect 756 69 768 87
rect 756 63 759 69
rect 765 63 768 69
rect 756 60 768 63
rect 804 93 816 96
rect 804 87 807 93
rect 813 87 816 93
rect 804 69 816 87
rect 804 63 807 69
rect 813 63 816 69
rect 804 60 816 63
rect 876 93 888 183
rect 876 87 879 93
rect 885 87 888 93
rect 876 69 888 87
rect 876 63 879 69
rect 885 63 888 69
rect 876 60 888 63
rect 924 93 936 96
rect 924 87 927 93
rect 933 87 936 93
rect 924 69 936 87
rect 924 63 927 69
rect 933 63 936 69
rect 924 60 936 63
rect 972 93 984 96
rect 972 87 975 93
rect 981 87 984 93
rect 972 69 984 87
rect 972 63 975 69
rect 981 63 984 69
rect 972 60 984 63
rect 1020 93 1032 96
rect 1020 87 1023 93
rect 1029 87 1032 93
rect 1020 69 1032 87
rect 1020 63 1023 69
rect 1029 63 1032 69
rect 1020 60 1032 63
rect 1092 93 1104 96
rect 1092 87 1095 93
rect 1101 87 1104 93
rect 1092 69 1104 87
rect 1092 63 1095 69
rect 1101 63 1104 69
rect 1092 60 1104 63
rect 1140 93 1152 96
rect 1140 87 1143 93
rect 1149 87 1152 93
rect 1140 69 1152 87
rect 1140 63 1143 69
rect 1149 63 1152 69
rect 1140 60 1152 63
rect 1188 93 1200 96
rect 1188 87 1191 93
rect 1197 87 1200 93
rect 1188 69 1200 87
rect 1188 63 1191 69
rect 1197 63 1200 69
rect 1188 60 1200 63
rect 1236 93 1248 96
rect 1236 87 1239 93
rect 1245 87 1248 93
rect 1236 69 1248 87
rect 1236 63 1239 69
rect 1245 63 1248 69
rect 1236 60 1248 63
<< labels >>
rlabel metal3 -24 408 -12 444 0 vdd
port 2 nsew
rlabel metal3 -24 12 -12 48 0 vss
port 3 nsew
rlabel metal3 -24 156 -12 168 0 x
rlabel metal3 -24 132 -12 144 0 y
rlabel metal3 -24 384 -12 396 0 bpa
rlabel metal3 -24 300 -12 312 0 bpb
rlabel metal3 -24 108 -12 120 0 bn0
rlabel metal3 -24 84 -12 96 0 bn
rlabel metal3 1272 204 1284 216 0 io
port 1 nsew
rlabel metal2 900 240 912 252 0 s
rlabel metal3 1272 228 1284 240 0 bnb
<< end >>
