magic
tech gf180mcuC
timestamp 1697453150
<< nwell >>
rect -90 486 1614 606
rect -90 342 1614 462
<< nmos >>
rect -48 12 -36 48
rect -24 12 -12 48
rect 0 12 12 48
rect 24 12 36 48
rect 48 12 60 48
rect 72 12 84 48
rect 96 12 108 48
rect 120 12 132 48
rect 144 12 156 48
rect 168 12 180 48
rect 192 12 204 48
rect 216 12 228 48
rect 240 12 252 48
rect 264 12 276 48
rect 288 12 300 48
rect 312 12 324 48
rect 336 12 348 48
rect 360 12 372 48
rect 384 12 396 48
rect 408 12 420 48
rect 432 12 444 48
rect 456 12 468 48
rect 480 12 492 48
rect 504 12 516 48
rect 528 12 540 48
rect 552 12 564 48
rect 576 12 588 48
rect 600 12 612 48
rect 624 12 636 48
rect 648 12 660 48
rect 672 12 684 48
rect 696 12 708 48
rect 720 12 732 48
rect 744 12 756 48
rect 768 12 780 48
rect 792 12 804 48
rect 816 12 828 48
rect 840 12 852 48
rect 864 12 876 48
rect 888 12 900 48
rect 912 12 924 48
rect 936 12 948 48
rect 960 12 972 48
rect 984 12 996 48
rect 1008 12 1020 48
rect 1032 12 1044 48
rect 1056 12 1068 48
rect 1080 12 1092 48
rect 1104 12 1116 48
rect 1128 12 1140 48
rect 1152 12 1164 48
rect 1176 12 1188 48
rect 1200 12 1212 48
rect 1224 12 1236 48
rect 1248 12 1260 48
rect 1272 12 1284 48
rect 1296 12 1308 48
rect 1320 12 1332 48
rect 1344 12 1356 48
rect 1368 12 1380 48
rect 1392 12 1404 48
rect 1416 12 1428 48
rect 1440 12 1452 48
rect 1464 12 1476 48
rect 1488 12 1500 48
rect 1512 12 1524 48
rect 1536 12 1548 48
rect 1560 12 1572 48
<< pmos >>
rect -48 396 -36 426
rect -24 396 -12 426
rect 0 396 12 426
rect 24 396 36 426
rect 48 396 60 426
rect 72 396 84 426
rect 96 396 108 426
rect 120 396 132 426
rect 144 396 156 426
rect 168 396 180 426
rect 192 396 204 426
rect 216 396 228 426
rect 240 396 252 426
rect 264 396 276 426
rect 288 396 300 426
rect 312 396 324 426
rect 336 396 348 426
rect 360 396 372 426
rect 384 396 396 426
rect 408 396 420 426
rect 432 396 444 426
rect 456 396 468 426
rect 480 396 492 426
rect 504 396 516 426
rect 528 396 540 426
rect 552 396 564 426
rect 576 396 588 426
rect 600 396 612 426
rect 624 396 636 426
rect 648 396 660 426
rect 672 396 684 426
rect 696 396 708 426
rect 720 396 732 426
rect 744 396 756 426
rect 768 396 780 426
rect 792 396 804 426
rect 816 396 828 426
rect 840 396 852 426
rect 864 396 876 426
rect 888 396 900 426
rect 912 396 924 426
rect 936 396 948 426
rect 960 396 972 426
rect 984 396 996 426
rect 1008 396 1020 426
rect 1032 396 1044 426
rect 1056 396 1068 426
rect 1080 396 1092 426
rect 1104 396 1116 426
rect 1128 396 1140 426
rect 1152 396 1164 426
rect 1176 396 1188 426
rect 1200 396 1212 426
rect 1224 396 1236 426
rect 1248 396 1260 426
rect 1272 396 1284 426
rect 1296 396 1308 426
rect 1320 396 1332 426
rect 1344 396 1356 426
rect 1368 396 1380 426
rect 1392 396 1404 426
rect 1416 396 1428 426
rect 1440 396 1452 426
rect 1464 396 1476 426
rect 1488 396 1500 426
rect 1512 396 1524 426
rect 1536 396 1548 426
rect 1560 396 1572 426
<< mvpmos >>
rect -48 516 -36 552
rect -24 516 -12 552
rect 0 516 12 552
rect 24 516 36 552
rect 48 516 60 552
rect 72 516 84 552
rect 96 516 108 552
rect 120 516 132 552
rect 144 516 156 552
rect 168 516 180 552
rect 192 516 204 552
rect 216 516 228 552
rect 240 516 252 552
rect 264 516 276 552
rect 288 516 300 552
rect 312 516 324 552
rect 336 516 348 552
rect 360 516 372 552
rect 384 516 396 552
rect 408 516 420 552
rect 432 516 444 552
rect 456 516 468 552
rect 480 516 492 552
rect 504 516 516 552
rect 528 516 540 552
rect 552 516 564 552
rect 576 516 588 552
rect 600 516 612 552
rect 624 516 636 552
rect 648 516 660 552
rect 672 516 684 552
rect 696 516 708 552
rect 720 516 732 552
rect 744 516 756 552
rect 768 516 780 552
rect 792 516 804 552
rect 816 516 828 552
rect 840 516 852 552
rect 864 516 876 552
rect 888 516 900 552
rect 912 516 924 552
rect 936 516 948 552
rect 960 516 972 552
rect 984 516 996 552
rect 1008 516 1020 552
rect 1032 516 1044 552
rect 1056 516 1068 552
rect 1080 516 1092 552
rect 1104 516 1116 552
rect 1128 516 1140 552
rect 1152 516 1164 552
rect 1176 516 1188 552
rect 1200 516 1212 552
rect 1224 516 1236 552
rect 1248 516 1260 552
rect 1272 516 1284 552
rect 1296 516 1308 552
rect 1320 516 1332 552
rect 1344 516 1356 552
rect 1368 516 1380 552
rect 1392 516 1404 552
rect 1416 516 1428 552
rect 1440 516 1452 552
rect 1464 516 1476 552
rect 1488 516 1500 552
rect 1512 516 1524 552
rect 1536 516 1548 552
rect 1560 516 1572 552
<< ndiff >>
rect -60 45 -48 48
rect -60 39 -57 45
rect -51 39 -48 45
rect -60 33 -48 39
rect -60 27 -57 33
rect -51 27 -48 33
rect -60 21 -48 27
rect -60 15 -57 21
rect -51 15 -48 21
rect -60 12 -48 15
rect -36 45 -24 48
rect -36 39 -33 45
rect -27 39 -24 45
rect -36 33 -24 39
rect -36 27 -33 33
rect -27 27 -24 33
rect -36 21 -24 27
rect -36 15 -33 21
rect -27 15 -24 21
rect -36 12 -24 15
rect -12 45 0 48
rect -12 39 -9 45
rect -3 39 0 45
rect -12 33 0 39
rect -12 27 -9 33
rect -3 27 0 33
rect -12 21 0 27
rect -12 15 -9 21
rect -3 15 0 21
rect -12 12 0 15
rect 12 12 24 48
rect 36 45 48 48
rect 36 39 39 45
rect 45 39 48 45
rect 36 33 48 39
rect 36 27 39 33
rect 45 27 48 33
rect 36 21 48 27
rect 36 15 39 21
rect 45 15 48 21
rect 36 12 48 15
rect 60 12 72 48
rect 84 45 96 48
rect 84 39 87 45
rect 93 39 96 45
rect 84 33 96 39
rect 84 27 87 33
rect 93 27 96 33
rect 84 21 96 27
rect 84 15 87 21
rect 93 15 96 21
rect 84 12 96 15
rect 108 12 120 48
rect 132 45 144 48
rect 132 39 135 45
rect 141 39 144 45
rect 132 33 144 39
rect 132 27 135 33
rect 141 27 144 33
rect 132 21 144 27
rect 132 15 135 21
rect 141 15 144 21
rect 132 12 144 15
rect 156 12 168 48
rect 180 45 192 48
rect 180 39 183 45
rect 189 39 192 45
rect 180 33 192 39
rect 180 27 183 33
rect 189 27 192 33
rect 180 21 192 27
rect 180 15 183 21
rect 189 15 192 21
rect 180 12 192 15
rect 204 12 216 48
rect 228 12 240 48
rect 252 12 264 48
rect 276 45 288 48
rect 276 39 279 45
rect 285 39 288 45
rect 276 33 288 39
rect 276 27 279 33
rect 285 27 288 33
rect 276 21 288 27
rect 276 15 279 21
rect 285 15 288 21
rect 276 12 288 15
rect 300 12 312 48
rect 324 12 336 48
rect 348 12 360 48
rect 372 45 384 48
rect 372 39 375 45
rect 381 39 384 45
rect 372 33 384 39
rect 372 27 375 33
rect 381 27 384 33
rect 372 21 384 27
rect 372 15 375 21
rect 381 15 384 21
rect 372 12 384 15
rect 396 12 408 48
rect 420 12 432 48
rect 444 12 456 48
rect 468 45 480 48
rect 468 39 471 45
rect 477 39 480 45
rect 468 33 480 39
rect 468 27 471 33
rect 477 27 480 33
rect 468 21 480 27
rect 468 15 471 21
rect 477 15 480 21
rect 468 12 480 15
rect 492 12 504 48
rect 516 12 528 48
rect 540 12 552 48
rect 564 45 576 48
rect 564 39 567 45
rect 573 39 576 45
rect 564 33 576 39
rect 564 27 567 33
rect 573 27 576 33
rect 564 21 576 27
rect 564 15 567 21
rect 573 15 576 21
rect 564 12 576 15
rect 588 12 600 48
rect 612 45 624 48
rect 612 39 615 45
rect 621 39 624 45
rect 612 33 624 39
rect 612 27 615 33
rect 621 27 624 33
rect 612 21 624 27
rect 612 15 615 21
rect 621 15 624 21
rect 612 12 624 15
rect 636 12 648 48
rect 660 45 672 48
rect 660 39 663 45
rect 669 39 672 45
rect 660 33 672 39
rect 660 27 663 33
rect 669 27 672 33
rect 660 21 672 27
rect 660 15 663 21
rect 669 15 672 21
rect 660 12 672 15
rect 684 12 696 48
rect 708 45 720 48
rect 708 39 711 45
rect 717 39 720 45
rect 708 33 720 39
rect 708 27 711 33
rect 717 27 720 33
rect 708 21 720 27
rect 708 15 711 21
rect 717 15 720 21
rect 708 12 720 15
rect 732 12 744 48
rect 756 45 768 48
rect 756 39 759 45
rect 765 39 768 45
rect 756 33 768 39
rect 756 27 759 33
rect 765 27 768 33
rect 756 21 768 27
rect 756 15 759 21
rect 765 15 768 21
rect 756 12 768 15
rect 780 12 792 48
rect 804 45 816 48
rect 804 39 807 45
rect 813 39 816 45
rect 804 33 816 39
rect 804 27 807 33
rect 813 27 816 33
rect 804 21 816 27
rect 804 15 807 21
rect 813 15 816 21
rect 804 12 816 15
rect 828 12 840 48
rect 852 45 864 48
rect 852 39 855 45
rect 861 39 864 45
rect 852 33 864 39
rect 852 27 855 33
rect 861 27 864 33
rect 852 21 864 27
rect 852 15 855 21
rect 861 15 864 21
rect 852 12 864 15
rect 876 12 888 48
rect 900 45 912 48
rect 900 39 903 45
rect 909 39 912 45
rect 900 33 912 39
rect 900 27 903 33
rect 909 27 912 33
rect 900 21 912 27
rect 900 15 903 21
rect 909 15 912 21
rect 900 12 912 15
rect 924 12 936 48
rect 948 45 960 48
rect 948 39 951 45
rect 957 39 960 45
rect 948 33 960 39
rect 948 27 951 33
rect 957 27 960 33
rect 948 21 960 27
rect 948 15 951 21
rect 957 15 960 21
rect 948 12 960 15
rect 972 12 984 48
rect 996 12 1008 48
rect 1020 12 1032 48
rect 1044 45 1056 48
rect 1044 39 1047 45
rect 1053 39 1056 45
rect 1044 33 1056 39
rect 1044 27 1047 33
rect 1053 27 1056 33
rect 1044 21 1056 27
rect 1044 15 1047 21
rect 1053 15 1056 21
rect 1044 12 1056 15
rect 1068 12 1080 48
rect 1092 12 1104 48
rect 1116 12 1128 48
rect 1140 45 1152 48
rect 1140 39 1143 45
rect 1149 39 1152 45
rect 1140 33 1152 39
rect 1140 27 1143 33
rect 1149 27 1152 33
rect 1140 21 1152 27
rect 1140 15 1143 21
rect 1149 15 1152 21
rect 1140 12 1152 15
rect 1164 12 1176 48
rect 1188 12 1200 48
rect 1212 12 1224 48
rect 1236 45 1248 48
rect 1236 39 1239 45
rect 1245 39 1248 45
rect 1236 33 1248 39
rect 1236 27 1239 33
rect 1245 27 1248 33
rect 1236 21 1248 27
rect 1236 15 1239 21
rect 1245 15 1248 21
rect 1236 12 1248 15
rect 1260 12 1272 48
rect 1284 12 1296 48
rect 1308 12 1320 48
rect 1332 45 1344 48
rect 1332 39 1335 45
rect 1341 39 1344 45
rect 1332 33 1344 39
rect 1332 27 1335 33
rect 1341 27 1344 33
rect 1332 21 1344 27
rect 1332 15 1335 21
rect 1341 15 1344 21
rect 1332 12 1344 15
rect 1356 12 1368 48
rect 1380 45 1392 48
rect 1380 39 1383 45
rect 1389 39 1392 45
rect 1380 33 1392 39
rect 1380 27 1383 33
rect 1389 27 1392 33
rect 1380 21 1392 27
rect 1380 15 1383 21
rect 1389 15 1392 21
rect 1380 12 1392 15
rect 1404 12 1416 48
rect 1428 45 1440 48
rect 1428 39 1431 45
rect 1437 39 1440 45
rect 1428 33 1440 39
rect 1428 27 1431 33
rect 1437 27 1440 33
rect 1428 21 1440 27
rect 1428 15 1431 21
rect 1437 15 1440 21
rect 1428 12 1440 15
rect 1452 12 1464 48
rect 1476 45 1488 48
rect 1476 39 1479 45
rect 1485 39 1488 45
rect 1476 33 1488 39
rect 1476 27 1479 33
rect 1485 27 1488 33
rect 1476 21 1488 27
rect 1476 15 1479 21
rect 1485 15 1488 21
rect 1476 12 1488 15
rect 1500 12 1512 48
rect 1524 45 1536 48
rect 1524 39 1527 45
rect 1533 39 1536 45
rect 1524 33 1536 39
rect 1524 27 1527 33
rect 1533 27 1536 33
rect 1524 21 1536 27
rect 1524 15 1527 21
rect 1533 15 1536 21
rect 1524 12 1536 15
rect 1548 45 1560 48
rect 1548 39 1551 45
rect 1557 39 1560 45
rect 1548 33 1560 39
rect 1548 27 1551 33
rect 1557 27 1560 33
rect 1548 21 1560 27
rect 1548 15 1551 21
rect 1557 15 1560 21
rect 1548 12 1560 15
rect 1572 45 1584 48
rect 1572 39 1575 45
rect 1581 39 1584 45
rect 1572 33 1584 39
rect 1572 27 1575 33
rect 1581 27 1584 33
rect 1572 21 1584 27
rect 1572 15 1575 21
rect 1581 15 1584 21
rect 1572 12 1584 15
<< pdiff >>
rect -60 417 -48 426
rect -60 411 -57 417
rect -51 411 -48 417
rect -60 405 -48 411
rect -60 399 -57 405
rect -51 399 -48 405
rect -60 396 -48 399
rect -36 417 -24 426
rect -36 411 -33 417
rect -27 411 -24 417
rect -36 405 -24 411
rect -36 399 -33 405
rect -27 399 -24 405
rect -36 396 -24 399
rect -12 417 0 426
rect -12 411 -9 417
rect -3 411 0 417
rect -12 405 0 411
rect -12 399 -9 405
rect -3 399 0 405
rect -12 396 0 399
rect 12 417 24 426
rect 12 411 15 417
rect 21 411 24 417
rect 12 405 24 411
rect 12 399 15 405
rect 21 399 24 405
rect 12 396 24 399
rect 36 417 48 426
rect 36 411 39 417
rect 45 411 48 417
rect 36 405 48 411
rect 36 399 39 405
rect 45 399 48 405
rect 36 396 48 399
rect 60 417 72 426
rect 60 411 63 417
rect 69 411 72 417
rect 60 405 72 411
rect 60 399 63 405
rect 69 399 72 405
rect 60 396 72 399
rect 84 417 96 426
rect 84 411 87 417
rect 93 411 96 417
rect 84 405 96 411
rect 84 399 87 405
rect 93 399 96 405
rect 84 396 96 399
rect 108 417 120 426
rect 108 411 111 417
rect 117 411 120 417
rect 108 405 120 411
rect 108 399 111 405
rect 117 399 120 405
rect 108 396 120 399
rect 132 417 144 426
rect 132 411 135 417
rect 141 411 144 417
rect 132 405 144 411
rect 132 399 135 405
rect 141 399 144 405
rect 132 396 144 399
rect 156 417 168 426
rect 156 411 159 417
rect 165 411 168 417
rect 156 405 168 411
rect 156 399 159 405
rect 165 399 168 405
rect 156 396 168 399
rect 180 417 192 426
rect 180 411 183 417
rect 189 411 192 417
rect 180 405 192 411
rect 180 399 183 405
rect 189 399 192 405
rect 180 396 192 399
rect 204 396 216 426
rect 228 417 240 426
rect 228 411 231 417
rect 237 411 240 417
rect 228 405 240 411
rect 228 399 231 405
rect 237 399 240 405
rect 228 396 240 399
rect 252 396 264 426
rect 276 417 288 426
rect 276 411 279 417
rect 285 411 288 417
rect 276 405 288 411
rect 276 399 279 405
rect 285 399 288 405
rect 276 396 288 399
rect 300 396 312 426
rect 324 417 336 426
rect 324 411 327 417
rect 333 411 336 417
rect 324 405 336 411
rect 324 399 327 405
rect 333 399 336 405
rect 324 396 336 399
rect 348 396 360 426
rect 372 417 384 426
rect 372 411 375 417
rect 381 411 384 417
rect 372 405 384 411
rect 372 399 375 405
rect 381 399 384 405
rect 372 396 384 399
rect 396 396 408 426
rect 420 417 432 426
rect 420 411 423 417
rect 429 411 432 417
rect 420 405 432 411
rect 420 399 423 405
rect 429 399 432 405
rect 420 396 432 399
rect 444 396 456 426
rect 468 417 480 426
rect 468 411 471 417
rect 477 411 480 417
rect 468 405 480 411
rect 468 399 471 405
rect 477 399 480 405
rect 468 396 480 399
rect 492 396 504 426
rect 516 417 528 426
rect 516 411 519 417
rect 525 411 528 417
rect 516 405 528 411
rect 516 399 519 405
rect 525 399 528 405
rect 516 396 528 399
rect 540 396 552 426
rect 564 417 576 426
rect 564 411 567 417
rect 573 411 576 417
rect 564 405 576 411
rect 564 399 567 405
rect 573 399 576 405
rect 564 396 576 399
rect 588 417 600 426
rect 588 411 591 417
rect 597 411 600 417
rect 588 405 600 411
rect 588 399 591 405
rect 597 399 600 405
rect 588 396 600 399
rect 612 417 624 426
rect 612 411 615 417
rect 621 411 624 417
rect 612 405 624 411
rect 612 399 615 405
rect 621 399 624 405
rect 612 396 624 399
rect 636 417 648 426
rect 636 411 639 417
rect 645 411 648 417
rect 636 405 648 411
rect 636 399 639 405
rect 645 399 648 405
rect 636 396 648 399
rect 660 417 672 426
rect 660 411 663 417
rect 669 411 672 417
rect 660 405 672 411
rect 660 399 663 405
rect 669 399 672 405
rect 660 396 672 399
rect 684 417 696 426
rect 684 411 687 417
rect 693 411 696 417
rect 684 405 696 411
rect 684 399 687 405
rect 693 399 696 405
rect 684 396 696 399
rect 708 417 720 426
rect 708 411 711 417
rect 717 411 720 417
rect 708 405 720 411
rect 708 399 711 405
rect 717 399 720 405
rect 708 396 720 399
rect 732 417 744 426
rect 732 411 735 417
rect 741 411 744 417
rect 732 405 744 411
rect 732 399 735 405
rect 741 399 744 405
rect 732 396 744 399
rect 756 417 768 426
rect 756 411 759 417
rect 765 411 768 417
rect 756 405 768 411
rect 756 399 759 405
rect 765 399 768 405
rect 756 396 768 399
rect 780 417 792 426
rect 780 411 783 417
rect 789 411 792 417
rect 780 405 792 411
rect 780 399 783 405
rect 789 399 792 405
rect 780 396 792 399
rect 804 417 816 426
rect 804 411 807 417
rect 813 411 816 417
rect 804 405 816 411
rect 804 399 807 405
rect 813 399 816 405
rect 804 396 816 399
rect 828 417 840 426
rect 828 411 831 417
rect 837 411 840 417
rect 828 405 840 411
rect 828 399 831 405
rect 837 399 840 405
rect 828 396 840 399
rect 852 417 864 426
rect 852 411 855 417
rect 861 411 864 417
rect 852 405 864 411
rect 852 399 855 405
rect 861 399 864 405
rect 852 396 864 399
rect 876 417 888 426
rect 876 411 879 417
rect 885 411 888 417
rect 876 405 888 411
rect 876 399 879 405
rect 885 399 888 405
rect 876 396 888 399
rect 900 417 912 426
rect 900 411 903 417
rect 909 411 912 417
rect 900 405 912 411
rect 900 399 903 405
rect 909 399 912 405
rect 900 396 912 399
rect 924 417 936 426
rect 924 411 927 417
rect 933 411 936 417
rect 924 405 936 411
rect 924 399 927 405
rect 933 399 936 405
rect 924 396 936 399
rect 948 417 960 426
rect 948 411 951 417
rect 957 411 960 417
rect 948 405 960 411
rect 948 399 951 405
rect 957 399 960 405
rect 948 396 960 399
rect 972 396 984 426
rect 996 417 1008 426
rect 996 411 999 417
rect 1005 411 1008 417
rect 996 405 1008 411
rect 996 399 999 405
rect 1005 399 1008 405
rect 996 396 1008 399
rect 1020 396 1032 426
rect 1044 417 1056 426
rect 1044 411 1047 417
rect 1053 411 1056 417
rect 1044 405 1056 411
rect 1044 399 1047 405
rect 1053 399 1056 405
rect 1044 396 1056 399
rect 1068 396 1080 426
rect 1092 417 1104 426
rect 1092 411 1095 417
rect 1101 411 1104 417
rect 1092 405 1104 411
rect 1092 399 1095 405
rect 1101 399 1104 405
rect 1092 396 1104 399
rect 1116 396 1128 426
rect 1140 417 1152 426
rect 1140 411 1143 417
rect 1149 411 1152 417
rect 1140 405 1152 411
rect 1140 399 1143 405
rect 1149 399 1152 405
rect 1140 396 1152 399
rect 1164 396 1176 426
rect 1188 417 1200 426
rect 1188 411 1191 417
rect 1197 411 1200 417
rect 1188 405 1200 411
rect 1188 399 1191 405
rect 1197 399 1200 405
rect 1188 396 1200 399
rect 1212 396 1224 426
rect 1236 417 1248 426
rect 1236 411 1239 417
rect 1245 411 1248 417
rect 1236 405 1248 411
rect 1236 399 1239 405
rect 1245 399 1248 405
rect 1236 396 1248 399
rect 1260 396 1272 426
rect 1284 417 1296 426
rect 1284 411 1287 417
rect 1293 411 1296 417
rect 1284 405 1296 411
rect 1284 399 1287 405
rect 1293 399 1296 405
rect 1284 396 1296 399
rect 1308 396 1320 426
rect 1332 417 1344 426
rect 1332 411 1335 417
rect 1341 411 1344 417
rect 1332 405 1344 411
rect 1332 399 1335 405
rect 1341 399 1344 405
rect 1332 396 1344 399
rect 1356 417 1368 426
rect 1356 411 1359 417
rect 1365 411 1368 417
rect 1356 405 1368 411
rect 1356 399 1359 405
rect 1365 399 1368 405
rect 1356 396 1368 399
rect 1380 417 1392 426
rect 1380 411 1383 417
rect 1389 411 1392 417
rect 1380 405 1392 411
rect 1380 399 1383 405
rect 1389 399 1392 405
rect 1380 396 1392 399
rect 1404 417 1416 426
rect 1404 411 1407 417
rect 1413 411 1416 417
rect 1404 405 1416 411
rect 1404 399 1407 405
rect 1413 399 1416 405
rect 1404 396 1416 399
rect 1428 417 1440 426
rect 1428 411 1431 417
rect 1437 411 1440 417
rect 1428 405 1440 411
rect 1428 399 1431 405
rect 1437 399 1440 405
rect 1428 396 1440 399
rect 1452 417 1464 426
rect 1452 411 1455 417
rect 1461 411 1464 417
rect 1452 405 1464 411
rect 1452 399 1455 405
rect 1461 399 1464 405
rect 1452 396 1464 399
rect 1476 417 1488 426
rect 1476 411 1479 417
rect 1485 411 1488 417
rect 1476 405 1488 411
rect 1476 399 1479 405
rect 1485 399 1488 405
rect 1476 396 1488 399
rect 1500 417 1512 426
rect 1500 411 1503 417
rect 1509 411 1512 417
rect 1500 405 1512 411
rect 1500 399 1503 405
rect 1509 399 1512 405
rect 1500 396 1512 399
rect 1524 417 1536 426
rect 1524 411 1527 417
rect 1533 411 1536 417
rect 1524 405 1536 411
rect 1524 399 1527 405
rect 1533 399 1536 405
rect 1524 396 1536 399
rect 1548 417 1560 426
rect 1548 411 1551 417
rect 1557 411 1560 417
rect 1548 405 1560 411
rect 1548 399 1551 405
rect 1557 399 1560 405
rect 1548 396 1560 399
rect 1572 417 1584 426
rect 1572 411 1575 417
rect 1581 411 1584 417
rect 1572 405 1584 411
rect 1572 399 1575 405
rect 1581 399 1584 405
rect 1572 396 1584 399
<< mvpdiff >>
rect -60 549 -48 552
rect -60 543 -57 549
rect -51 543 -48 549
rect -60 537 -48 543
rect -60 531 -57 537
rect -51 531 -48 537
rect -60 525 -48 531
rect -60 519 -57 525
rect -51 519 -48 525
rect -60 516 -48 519
rect -36 549 -24 552
rect -36 543 -33 549
rect -27 543 -24 549
rect -36 537 -24 543
rect -36 531 -33 537
rect -27 531 -24 537
rect -36 525 -24 531
rect -36 519 -33 525
rect -27 519 -24 525
rect -36 516 -24 519
rect -12 549 0 552
rect -12 543 -9 549
rect -3 543 0 549
rect -12 537 0 543
rect -12 531 -9 537
rect -3 531 0 537
rect -12 525 0 531
rect -12 519 -9 525
rect -3 519 0 525
rect -12 516 0 519
rect 12 549 24 552
rect 12 543 15 549
rect 21 543 24 549
rect 12 537 24 543
rect 12 531 15 537
rect 21 531 24 537
rect 12 525 24 531
rect 12 519 15 525
rect 21 519 24 525
rect 12 516 24 519
rect 36 549 48 552
rect 36 543 39 549
rect 45 543 48 549
rect 36 537 48 543
rect 36 531 39 537
rect 45 531 48 537
rect 36 525 48 531
rect 36 519 39 525
rect 45 519 48 525
rect 36 516 48 519
rect 60 549 72 552
rect 60 543 63 549
rect 69 543 72 549
rect 60 537 72 543
rect 60 531 63 537
rect 69 531 72 537
rect 60 525 72 531
rect 60 519 63 525
rect 69 519 72 525
rect 60 516 72 519
rect 84 549 96 552
rect 84 543 87 549
rect 93 543 96 549
rect 84 537 96 543
rect 84 531 87 537
rect 93 531 96 537
rect 84 525 96 531
rect 84 519 87 525
rect 93 519 96 525
rect 84 516 96 519
rect 108 549 120 552
rect 108 543 111 549
rect 117 543 120 549
rect 108 537 120 543
rect 108 531 111 537
rect 117 531 120 537
rect 108 525 120 531
rect 108 519 111 525
rect 117 519 120 525
rect 108 516 120 519
rect 132 549 144 552
rect 132 543 135 549
rect 141 543 144 549
rect 132 537 144 543
rect 132 531 135 537
rect 141 531 144 537
rect 132 525 144 531
rect 132 519 135 525
rect 141 519 144 525
rect 132 516 144 519
rect 156 549 168 552
rect 156 543 159 549
rect 165 543 168 549
rect 156 537 168 543
rect 156 531 159 537
rect 165 531 168 537
rect 156 525 168 531
rect 156 519 159 525
rect 165 519 168 525
rect 156 516 168 519
rect 180 549 192 552
rect 180 543 183 549
rect 189 543 192 549
rect 180 537 192 543
rect 180 531 183 537
rect 189 531 192 537
rect 180 525 192 531
rect 180 519 183 525
rect 189 519 192 525
rect 180 516 192 519
rect 204 549 216 552
rect 204 543 207 549
rect 213 543 216 549
rect 204 537 216 543
rect 204 531 207 537
rect 213 531 216 537
rect 204 525 216 531
rect 204 519 207 525
rect 213 519 216 525
rect 204 516 216 519
rect 228 549 240 552
rect 228 543 231 549
rect 237 543 240 549
rect 228 537 240 543
rect 228 531 231 537
rect 237 531 240 537
rect 228 525 240 531
rect 228 519 231 525
rect 237 519 240 525
rect 228 516 240 519
rect 252 549 264 552
rect 252 543 255 549
rect 261 543 264 549
rect 252 537 264 543
rect 252 531 255 537
rect 261 531 264 537
rect 252 525 264 531
rect 252 519 255 525
rect 261 519 264 525
rect 252 516 264 519
rect 276 549 288 552
rect 276 543 279 549
rect 285 543 288 549
rect 276 537 288 543
rect 276 531 279 537
rect 285 531 288 537
rect 276 525 288 531
rect 276 519 279 525
rect 285 519 288 525
rect 276 516 288 519
rect 300 549 312 552
rect 300 543 303 549
rect 309 543 312 549
rect 300 537 312 543
rect 300 531 303 537
rect 309 531 312 537
rect 300 525 312 531
rect 300 519 303 525
rect 309 519 312 525
rect 300 516 312 519
rect 324 549 336 552
rect 324 543 327 549
rect 333 543 336 549
rect 324 537 336 543
rect 324 531 327 537
rect 333 531 336 537
rect 324 525 336 531
rect 324 519 327 525
rect 333 519 336 525
rect 324 516 336 519
rect 348 549 360 552
rect 348 543 351 549
rect 357 543 360 549
rect 348 537 360 543
rect 348 531 351 537
rect 357 531 360 537
rect 348 525 360 531
rect 348 519 351 525
rect 357 519 360 525
rect 348 516 360 519
rect 372 549 384 552
rect 372 543 375 549
rect 381 543 384 549
rect 372 537 384 543
rect 372 531 375 537
rect 381 531 384 537
rect 372 525 384 531
rect 372 519 375 525
rect 381 519 384 525
rect 372 516 384 519
rect 396 549 408 552
rect 396 543 399 549
rect 405 543 408 549
rect 396 537 408 543
rect 396 531 399 537
rect 405 531 408 537
rect 396 525 408 531
rect 396 519 399 525
rect 405 519 408 525
rect 396 516 408 519
rect 420 549 432 552
rect 420 543 423 549
rect 429 543 432 549
rect 420 537 432 543
rect 420 531 423 537
rect 429 531 432 537
rect 420 525 432 531
rect 420 519 423 525
rect 429 519 432 525
rect 420 516 432 519
rect 444 549 456 552
rect 444 543 447 549
rect 453 543 456 549
rect 444 537 456 543
rect 444 531 447 537
rect 453 531 456 537
rect 444 525 456 531
rect 444 519 447 525
rect 453 519 456 525
rect 444 516 456 519
rect 468 549 480 552
rect 468 543 471 549
rect 477 543 480 549
rect 468 537 480 543
rect 468 531 471 537
rect 477 531 480 537
rect 468 525 480 531
rect 468 519 471 525
rect 477 519 480 525
rect 468 516 480 519
rect 492 549 504 552
rect 492 543 495 549
rect 501 543 504 549
rect 492 537 504 543
rect 492 531 495 537
rect 501 531 504 537
rect 492 525 504 531
rect 492 519 495 525
rect 501 519 504 525
rect 492 516 504 519
rect 516 549 528 552
rect 516 543 519 549
rect 525 543 528 549
rect 516 537 528 543
rect 516 531 519 537
rect 525 531 528 537
rect 516 525 528 531
rect 516 519 519 525
rect 525 519 528 525
rect 516 516 528 519
rect 540 549 552 552
rect 540 543 543 549
rect 549 543 552 549
rect 540 537 552 543
rect 540 531 543 537
rect 549 531 552 537
rect 540 525 552 531
rect 540 519 543 525
rect 549 519 552 525
rect 540 516 552 519
rect 564 549 576 552
rect 564 543 567 549
rect 573 543 576 549
rect 564 537 576 543
rect 564 531 567 537
rect 573 531 576 537
rect 564 525 576 531
rect 564 519 567 525
rect 573 519 576 525
rect 564 516 576 519
rect 588 549 600 552
rect 588 543 591 549
rect 597 543 600 549
rect 588 537 600 543
rect 588 531 591 537
rect 597 531 600 537
rect 588 525 600 531
rect 588 519 591 525
rect 597 519 600 525
rect 588 516 600 519
rect 612 549 624 552
rect 612 543 615 549
rect 621 543 624 549
rect 612 537 624 543
rect 612 531 615 537
rect 621 531 624 537
rect 612 525 624 531
rect 612 519 615 525
rect 621 519 624 525
rect 612 516 624 519
rect 636 549 648 552
rect 636 543 639 549
rect 645 543 648 549
rect 636 537 648 543
rect 636 531 639 537
rect 645 531 648 537
rect 636 525 648 531
rect 636 519 639 525
rect 645 519 648 525
rect 636 516 648 519
rect 660 549 672 552
rect 660 543 663 549
rect 669 543 672 549
rect 660 537 672 543
rect 660 531 663 537
rect 669 531 672 537
rect 660 525 672 531
rect 660 519 663 525
rect 669 519 672 525
rect 660 516 672 519
rect 684 549 696 552
rect 684 543 687 549
rect 693 543 696 549
rect 684 537 696 543
rect 684 531 687 537
rect 693 531 696 537
rect 684 525 696 531
rect 684 519 687 525
rect 693 519 696 525
rect 684 516 696 519
rect 708 549 720 552
rect 708 543 711 549
rect 717 543 720 549
rect 708 537 720 543
rect 708 531 711 537
rect 717 531 720 537
rect 708 525 720 531
rect 708 519 711 525
rect 717 519 720 525
rect 708 516 720 519
rect 732 549 744 552
rect 732 543 735 549
rect 741 543 744 549
rect 732 537 744 543
rect 732 531 735 537
rect 741 531 744 537
rect 732 525 744 531
rect 732 519 735 525
rect 741 519 744 525
rect 732 516 744 519
rect 756 549 768 552
rect 756 543 759 549
rect 765 543 768 549
rect 756 537 768 543
rect 756 531 759 537
rect 765 531 768 537
rect 756 525 768 531
rect 756 519 759 525
rect 765 519 768 525
rect 756 516 768 519
rect 780 549 792 552
rect 780 543 783 549
rect 789 543 792 549
rect 780 537 792 543
rect 780 531 783 537
rect 789 531 792 537
rect 780 525 792 531
rect 780 519 783 525
rect 789 519 792 525
rect 780 516 792 519
rect 804 549 816 552
rect 804 543 807 549
rect 813 543 816 549
rect 804 537 816 543
rect 804 531 807 537
rect 813 531 816 537
rect 804 525 816 531
rect 804 519 807 525
rect 813 519 816 525
rect 804 516 816 519
rect 828 549 840 552
rect 828 543 831 549
rect 837 543 840 549
rect 828 537 840 543
rect 828 531 831 537
rect 837 531 840 537
rect 828 525 840 531
rect 828 519 831 525
rect 837 519 840 525
rect 828 516 840 519
rect 852 549 864 552
rect 852 543 855 549
rect 861 543 864 549
rect 852 537 864 543
rect 852 531 855 537
rect 861 531 864 537
rect 852 525 864 531
rect 852 519 855 525
rect 861 519 864 525
rect 852 516 864 519
rect 876 549 888 552
rect 876 543 879 549
rect 885 543 888 549
rect 876 537 888 543
rect 876 531 879 537
rect 885 531 888 537
rect 876 525 888 531
rect 876 519 879 525
rect 885 519 888 525
rect 876 516 888 519
rect 900 549 912 552
rect 900 543 903 549
rect 909 543 912 549
rect 900 537 912 543
rect 900 531 903 537
rect 909 531 912 537
rect 900 525 912 531
rect 900 519 903 525
rect 909 519 912 525
rect 900 516 912 519
rect 924 549 936 552
rect 924 543 927 549
rect 933 543 936 549
rect 924 537 936 543
rect 924 531 927 537
rect 933 531 936 537
rect 924 525 936 531
rect 924 519 927 525
rect 933 519 936 525
rect 924 516 936 519
rect 948 549 960 552
rect 948 543 951 549
rect 957 543 960 549
rect 948 537 960 543
rect 948 531 951 537
rect 957 531 960 537
rect 948 525 960 531
rect 948 519 951 525
rect 957 519 960 525
rect 948 516 960 519
rect 972 549 984 552
rect 972 543 975 549
rect 981 543 984 549
rect 972 537 984 543
rect 972 531 975 537
rect 981 531 984 537
rect 972 525 984 531
rect 972 519 975 525
rect 981 519 984 525
rect 972 516 984 519
rect 996 549 1008 552
rect 996 543 999 549
rect 1005 543 1008 549
rect 996 537 1008 543
rect 996 531 999 537
rect 1005 531 1008 537
rect 996 525 1008 531
rect 996 519 999 525
rect 1005 519 1008 525
rect 996 516 1008 519
rect 1020 549 1032 552
rect 1020 543 1023 549
rect 1029 543 1032 549
rect 1020 537 1032 543
rect 1020 531 1023 537
rect 1029 531 1032 537
rect 1020 525 1032 531
rect 1020 519 1023 525
rect 1029 519 1032 525
rect 1020 516 1032 519
rect 1044 549 1056 552
rect 1044 543 1047 549
rect 1053 543 1056 549
rect 1044 537 1056 543
rect 1044 531 1047 537
rect 1053 531 1056 537
rect 1044 525 1056 531
rect 1044 519 1047 525
rect 1053 519 1056 525
rect 1044 516 1056 519
rect 1068 549 1080 552
rect 1068 543 1071 549
rect 1077 543 1080 549
rect 1068 537 1080 543
rect 1068 531 1071 537
rect 1077 531 1080 537
rect 1068 525 1080 531
rect 1068 519 1071 525
rect 1077 519 1080 525
rect 1068 516 1080 519
rect 1092 549 1104 552
rect 1092 543 1095 549
rect 1101 543 1104 549
rect 1092 537 1104 543
rect 1092 531 1095 537
rect 1101 531 1104 537
rect 1092 525 1104 531
rect 1092 519 1095 525
rect 1101 519 1104 525
rect 1092 516 1104 519
rect 1116 549 1128 552
rect 1116 543 1119 549
rect 1125 543 1128 549
rect 1116 537 1128 543
rect 1116 531 1119 537
rect 1125 531 1128 537
rect 1116 525 1128 531
rect 1116 519 1119 525
rect 1125 519 1128 525
rect 1116 516 1128 519
rect 1140 549 1152 552
rect 1140 543 1143 549
rect 1149 543 1152 549
rect 1140 537 1152 543
rect 1140 531 1143 537
rect 1149 531 1152 537
rect 1140 525 1152 531
rect 1140 519 1143 525
rect 1149 519 1152 525
rect 1140 516 1152 519
rect 1164 549 1176 552
rect 1164 543 1167 549
rect 1173 543 1176 549
rect 1164 537 1176 543
rect 1164 531 1167 537
rect 1173 531 1176 537
rect 1164 525 1176 531
rect 1164 519 1167 525
rect 1173 519 1176 525
rect 1164 516 1176 519
rect 1188 549 1200 552
rect 1188 543 1191 549
rect 1197 543 1200 549
rect 1188 537 1200 543
rect 1188 531 1191 537
rect 1197 531 1200 537
rect 1188 525 1200 531
rect 1188 519 1191 525
rect 1197 519 1200 525
rect 1188 516 1200 519
rect 1212 549 1224 552
rect 1212 543 1215 549
rect 1221 543 1224 549
rect 1212 537 1224 543
rect 1212 531 1215 537
rect 1221 531 1224 537
rect 1212 525 1224 531
rect 1212 519 1215 525
rect 1221 519 1224 525
rect 1212 516 1224 519
rect 1236 549 1248 552
rect 1236 543 1239 549
rect 1245 543 1248 549
rect 1236 537 1248 543
rect 1236 531 1239 537
rect 1245 531 1248 537
rect 1236 525 1248 531
rect 1236 519 1239 525
rect 1245 519 1248 525
rect 1236 516 1248 519
rect 1260 549 1272 552
rect 1260 543 1263 549
rect 1269 543 1272 549
rect 1260 537 1272 543
rect 1260 531 1263 537
rect 1269 531 1272 537
rect 1260 525 1272 531
rect 1260 519 1263 525
rect 1269 519 1272 525
rect 1260 516 1272 519
rect 1284 549 1296 552
rect 1284 543 1287 549
rect 1293 543 1296 549
rect 1284 537 1296 543
rect 1284 531 1287 537
rect 1293 531 1296 537
rect 1284 525 1296 531
rect 1284 519 1287 525
rect 1293 519 1296 525
rect 1284 516 1296 519
rect 1308 549 1320 552
rect 1308 543 1311 549
rect 1317 543 1320 549
rect 1308 537 1320 543
rect 1308 531 1311 537
rect 1317 531 1320 537
rect 1308 525 1320 531
rect 1308 519 1311 525
rect 1317 519 1320 525
rect 1308 516 1320 519
rect 1332 549 1344 552
rect 1332 543 1335 549
rect 1341 543 1344 549
rect 1332 537 1344 543
rect 1332 531 1335 537
rect 1341 531 1344 537
rect 1332 525 1344 531
rect 1332 519 1335 525
rect 1341 519 1344 525
rect 1332 516 1344 519
rect 1356 549 1368 552
rect 1356 543 1359 549
rect 1365 543 1368 549
rect 1356 537 1368 543
rect 1356 531 1359 537
rect 1365 531 1368 537
rect 1356 525 1368 531
rect 1356 519 1359 525
rect 1365 519 1368 525
rect 1356 516 1368 519
rect 1380 549 1392 552
rect 1380 543 1383 549
rect 1389 543 1392 549
rect 1380 537 1392 543
rect 1380 531 1383 537
rect 1389 531 1392 537
rect 1380 525 1392 531
rect 1380 519 1383 525
rect 1389 519 1392 525
rect 1380 516 1392 519
rect 1404 549 1416 552
rect 1404 543 1407 549
rect 1413 543 1416 549
rect 1404 537 1416 543
rect 1404 531 1407 537
rect 1413 531 1416 537
rect 1404 525 1416 531
rect 1404 519 1407 525
rect 1413 519 1416 525
rect 1404 516 1416 519
rect 1428 549 1440 552
rect 1428 543 1431 549
rect 1437 543 1440 549
rect 1428 537 1440 543
rect 1428 531 1431 537
rect 1437 531 1440 537
rect 1428 525 1440 531
rect 1428 519 1431 525
rect 1437 519 1440 525
rect 1428 516 1440 519
rect 1452 549 1464 552
rect 1452 543 1455 549
rect 1461 543 1464 549
rect 1452 537 1464 543
rect 1452 531 1455 537
rect 1461 531 1464 537
rect 1452 525 1464 531
rect 1452 519 1455 525
rect 1461 519 1464 525
rect 1452 516 1464 519
rect 1476 549 1488 552
rect 1476 543 1479 549
rect 1485 543 1488 549
rect 1476 537 1488 543
rect 1476 531 1479 537
rect 1485 531 1488 537
rect 1476 525 1488 531
rect 1476 519 1479 525
rect 1485 519 1488 525
rect 1476 516 1488 519
rect 1500 549 1512 552
rect 1500 543 1503 549
rect 1509 543 1512 549
rect 1500 537 1512 543
rect 1500 531 1503 537
rect 1509 531 1512 537
rect 1500 525 1512 531
rect 1500 519 1503 525
rect 1509 519 1512 525
rect 1500 516 1512 519
rect 1524 549 1536 552
rect 1524 543 1527 549
rect 1533 543 1536 549
rect 1524 537 1536 543
rect 1524 531 1527 537
rect 1533 531 1536 537
rect 1524 525 1536 531
rect 1524 519 1527 525
rect 1533 519 1536 525
rect 1524 516 1536 519
rect 1548 549 1560 552
rect 1548 543 1551 549
rect 1557 543 1560 549
rect 1548 537 1560 543
rect 1548 531 1551 537
rect 1557 531 1560 537
rect 1548 525 1560 531
rect 1548 519 1551 525
rect 1557 519 1560 525
rect 1548 516 1560 519
rect 1572 549 1584 552
rect 1572 543 1575 549
rect 1581 543 1584 549
rect 1572 537 1584 543
rect 1572 531 1575 537
rect 1581 531 1584 537
rect 1572 525 1584 531
rect 1572 519 1575 525
rect 1581 519 1584 525
rect 1572 516 1584 519
<< ndiffc >>
rect -57 39 -51 45
rect -57 27 -51 33
rect -57 15 -51 21
rect -33 39 -27 45
rect -33 27 -27 33
rect -33 15 -27 21
rect -9 39 -3 45
rect -9 27 -3 33
rect -9 15 -3 21
rect 39 39 45 45
rect 39 27 45 33
rect 39 15 45 21
rect 87 39 93 45
rect 87 27 93 33
rect 87 15 93 21
rect 135 39 141 45
rect 135 27 141 33
rect 135 15 141 21
rect 183 39 189 45
rect 183 27 189 33
rect 183 15 189 21
rect 279 39 285 45
rect 279 27 285 33
rect 279 15 285 21
rect 375 39 381 45
rect 375 27 381 33
rect 375 15 381 21
rect 471 39 477 45
rect 471 27 477 33
rect 471 15 477 21
rect 567 39 573 45
rect 567 27 573 33
rect 567 15 573 21
rect 615 39 621 45
rect 615 27 621 33
rect 615 15 621 21
rect 663 39 669 45
rect 663 27 669 33
rect 663 15 669 21
rect 711 39 717 45
rect 711 27 717 33
rect 711 15 717 21
rect 759 39 765 45
rect 759 27 765 33
rect 759 15 765 21
rect 807 39 813 45
rect 807 27 813 33
rect 807 15 813 21
rect 855 39 861 45
rect 855 27 861 33
rect 855 15 861 21
rect 903 39 909 45
rect 903 27 909 33
rect 903 15 909 21
rect 951 39 957 45
rect 951 27 957 33
rect 951 15 957 21
rect 1047 39 1053 45
rect 1047 27 1053 33
rect 1047 15 1053 21
rect 1143 39 1149 45
rect 1143 27 1149 33
rect 1143 15 1149 21
rect 1239 39 1245 45
rect 1239 27 1245 33
rect 1239 15 1245 21
rect 1335 39 1341 45
rect 1335 27 1341 33
rect 1335 15 1341 21
rect 1383 39 1389 45
rect 1383 27 1389 33
rect 1383 15 1389 21
rect 1431 39 1437 45
rect 1431 27 1437 33
rect 1431 15 1437 21
rect 1479 39 1485 45
rect 1479 27 1485 33
rect 1479 15 1485 21
rect 1527 39 1533 45
rect 1527 27 1533 33
rect 1527 15 1533 21
rect 1551 39 1557 45
rect 1551 27 1557 33
rect 1551 15 1557 21
rect 1575 39 1581 45
rect 1575 27 1581 33
rect 1575 15 1581 21
<< pdiffc >>
rect -57 411 -51 417
rect -57 399 -51 405
rect -33 411 -27 417
rect -33 399 -27 405
rect -9 411 -3 417
rect -9 399 -3 405
rect 15 411 21 417
rect 15 399 21 405
rect 39 411 45 417
rect 39 399 45 405
rect 63 411 69 417
rect 63 399 69 405
rect 87 411 93 417
rect 87 399 93 405
rect 111 411 117 417
rect 111 399 117 405
rect 135 411 141 417
rect 135 399 141 405
rect 159 411 165 417
rect 159 399 165 405
rect 183 411 189 417
rect 183 399 189 405
rect 231 411 237 417
rect 231 399 237 405
rect 279 411 285 417
rect 279 399 285 405
rect 327 411 333 417
rect 327 399 333 405
rect 375 411 381 417
rect 375 399 381 405
rect 423 411 429 417
rect 423 399 429 405
rect 471 411 477 417
rect 471 399 477 405
rect 519 411 525 417
rect 519 399 525 405
rect 567 411 573 417
rect 567 399 573 405
rect 591 411 597 417
rect 591 399 597 405
rect 615 411 621 417
rect 615 399 621 405
rect 639 411 645 417
rect 639 399 645 405
rect 663 411 669 417
rect 663 399 669 405
rect 687 411 693 417
rect 687 399 693 405
rect 711 411 717 417
rect 711 399 717 405
rect 735 411 741 417
rect 735 399 741 405
rect 759 411 765 417
rect 759 399 765 405
rect 783 411 789 417
rect 783 399 789 405
rect 807 411 813 417
rect 807 399 813 405
rect 831 411 837 417
rect 831 399 837 405
rect 855 411 861 417
rect 855 399 861 405
rect 879 411 885 417
rect 879 399 885 405
rect 903 411 909 417
rect 903 399 909 405
rect 927 411 933 417
rect 927 399 933 405
rect 951 411 957 417
rect 951 399 957 405
rect 999 411 1005 417
rect 999 399 1005 405
rect 1047 411 1053 417
rect 1047 399 1053 405
rect 1095 411 1101 417
rect 1095 399 1101 405
rect 1143 411 1149 417
rect 1143 399 1149 405
rect 1191 411 1197 417
rect 1191 399 1197 405
rect 1239 411 1245 417
rect 1239 399 1245 405
rect 1287 411 1293 417
rect 1287 399 1293 405
rect 1335 411 1341 417
rect 1335 399 1341 405
rect 1359 411 1365 417
rect 1359 399 1365 405
rect 1383 411 1389 417
rect 1383 399 1389 405
rect 1407 411 1413 417
rect 1407 399 1413 405
rect 1431 411 1437 417
rect 1431 399 1437 405
rect 1455 411 1461 417
rect 1455 399 1461 405
rect 1479 411 1485 417
rect 1479 399 1485 405
rect 1503 411 1509 417
rect 1503 399 1509 405
rect 1527 411 1533 417
rect 1527 399 1533 405
rect 1551 411 1557 417
rect 1551 399 1557 405
rect 1575 411 1581 417
rect 1575 399 1581 405
<< mvpdiffc >>
rect -57 543 -51 549
rect -57 531 -51 537
rect -57 519 -51 525
rect -33 543 -27 549
rect -33 531 -27 537
rect -33 519 -27 525
rect -9 543 -3 549
rect -9 531 -3 537
rect -9 519 -3 525
rect 15 543 21 549
rect 15 531 21 537
rect 15 519 21 525
rect 39 543 45 549
rect 39 531 45 537
rect 39 519 45 525
rect 63 543 69 549
rect 63 531 69 537
rect 63 519 69 525
rect 87 543 93 549
rect 87 531 93 537
rect 87 519 93 525
rect 111 543 117 549
rect 111 531 117 537
rect 111 519 117 525
rect 135 543 141 549
rect 135 531 141 537
rect 135 519 141 525
rect 159 543 165 549
rect 159 531 165 537
rect 159 519 165 525
rect 183 543 189 549
rect 183 531 189 537
rect 183 519 189 525
rect 207 543 213 549
rect 207 531 213 537
rect 207 519 213 525
rect 231 543 237 549
rect 231 531 237 537
rect 231 519 237 525
rect 255 543 261 549
rect 255 531 261 537
rect 255 519 261 525
rect 279 543 285 549
rect 279 531 285 537
rect 279 519 285 525
rect 303 543 309 549
rect 303 531 309 537
rect 303 519 309 525
rect 327 543 333 549
rect 327 531 333 537
rect 327 519 333 525
rect 351 543 357 549
rect 351 531 357 537
rect 351 519 357 525
rect 375 543 381 549
rect 375 531 381 537
rect 375 519 381 525
rect 399 543 405 549
rect 399 531 405 537
rect 399 519 405 525
rect 423 543 429 549
rect 423 531 429 537
rect 423 519 429 525
rect 447 543 453 549
rect 447 531 453 537
rect 447 519 453 525
rect 471 543 477 549
rect 471 531 477 537
rect 471 519 477 525
rect 495 543 501 549
rect 495 531 501 537
rect 495 519 501 525
rect 519 543 525 549
rect 519 531 525 537
rect 519 519 525 525
rect 543 543 549 549
rect 543 531 549 537
rect 543 519 549 525
rect 567 543 573 549
rect 567 531 573 537
rect 567 519 573 525
rect 591 543 597 549
rect 591 531 597 537
rect 591 519 597 525
rect 615 543 621 549
rect 615 531 621 537
rect 615 519 621 525
rect 639 543 645 549
rect 639 531 645 537
rect 639 519 645 525
rect 663 543 669 549
rect 663 531 669 537
rect 663 519 669 525
rect 687 543 693 549
rect 687 531 693 537
rect 687 519 693 525
rect 711 543 717 549
rect 711 531 717 537
rect 711 519 717 525
rect 735 543 741 549
rect 735 531 741 537
rect 735 519 741 525
rect 759 543 765 549
rect 759 531 765 537
rect 759 519 765 525
rect 783 543 789 549
rect 783 531 789 537
rect 783 519 789 525
rect 807 543 813 549
rect 807 531 813 537
rect 807 519 813 525
rect 831 543 837 549
rect 831 531 837 537
rect 831 519 837 525
rect 855 543 861 549
rect 855 531 861 537
rect 855 519 861 525
rect 879 543 885 549
rect 879 531 885 537
rect 879 519 885 525
rect 903 543 909 549
rect 903 531 909 537
rect 903 519 909 525
rect 927 543 933 549
rect 927 531 933 537
rect 927 519 933 525
rect 951 543 957 549
rect 951 531 957 537
rect 951 519 957 525
rect 975 543 981 549
rect 975 531 981 537
rect 975 519 981 525
rect 999 543 1005 549
rect 999 531 1005 537
rect 999 519 1005 525
rect 1023 543 1029 549
rect 1023 531 1029 537
rect 1023 519 1029 525
rect 1047 543 1053 549
rect 1047 531 1053 537
rect 1047 519 1053 525
rect 1071 543 1077 549
rect 1071 531 1077 537
rect 1071 519 1077 525
rect 1095 543 1101 549
rect 1095 531 1101 537
rect 1095 519 1101 525
rect 1119 543 1125 549
rect 1119 531 1125 537
rect 1119 519 1125 525
rect 1143 543 1149 549
rect 1143 531 1149 537
rect 1143 519 1149 525
rect 1167 543 1173 549
rect 1167 531 1173 537
rect 1167 519 1173 525
rect 1191 543 1197 549
rect 1191 531 1197 537
rect 1191 519 1197 525
rect 1215 543 1221 549
rect 1215 531 1221 537
rect 1215 519 1221 525
rect 1239 543 1245 549
rect 1239 531 1245 537
rect 1239 519 1245 525
rect 1263 543 1269 549
rect 1263 531 1269 537
rect 1263 519 1269 525
rect 1287 543 1293 549
rect 1287 531 1293 537
rect 1287 519 1293 525
rect 1311 543 1317 549
rect 1311 531 1317 537
rect 1311 519 1317 525
rect 1335 543 1341 549
rect 1335 531 1341 537
rect 1335 519 1341 525
rect 1359 543 1365 549
rect 1359 531 1365 537
rect 1359 519 1365 525
rect 1383 543 1389 549
rect 1383 531 1389 537
rect 1383 519 1389 525
rect 1407 543 1413 549
rect 1407 531 1413 537
rect 1407 519 1413 525
rect 1431 543 1437 549
rect 1431 531 1437 537
rect 1431 519 1437 525
rect 1455 543 1461 549
rect 1455 531 1461 537
rect 1455 519 1461 525
rect 1479 543 1485 549
rect 1479 531 1485 537
rect 1479 519 1485 525
rect 1503 543 1509 549
rect 1503 531 1509 537
rect 1503 519 1509 525
rect 1527 543 1533 549
rect 1527 531 1533 537
rect 1527 519 1533 525
rect 1551 543 1557 549
rect 1551 531 1557 537
rect 1551 519 1557 525
rect 1575 543 1581 549
rect 1575 531 1581 537
rect 1575 519 1581 525
<< psubdiff >>
rect -108 621 1632 624
rect -108 615 -105 621
rect -99 615 -93 621
rect -87 615 -81 621
rect -75 615 -69 621
rect -63 615 -57 621
rect -51 615 -45 621
rect -39 615 -33 621
rect -27 615 -21 621
rect -15 615 -9 621
rect -3 615 3 621
rect 9 615 15 621
rect 21 615 27 621
rect 33 615 39 621
rect 45 615 51 621
rect 57 615 63 621
rect 69 615 75 621
rect 81 615 87 621
rect 93 615 99 621
rect 105 615 111 621
rect 117 615 123 621
rect 129 615 135 621
rect 141 615 147 621
rect 153 615 159 621
rect 165 615 171 621
rect 177 615 183 621
rect 189 615 195 621
rect 201 615 207 621
rect 213 615 219 621
rect 225 615 231 621
rect 237 615 243 621
rect 249 615 255 621
rect 261 615 267 621
rect 273 615 279 621
rect 285 615 291 621
rect 297 615 303 621
rect 309 615 315 621
rect 321 615 327 621
rect 333 615 339 621
rect 345 615 351 621
rect 357 615 363 621
rect 369 615 375 621
rect 381 615 387 621
rect 393 615 399 621
rect 405 615 411 621
rect 417 615 423 621
rect 429 615 435 621
rect 441 615 447 621
rect 453 615 459 621
rect 465 615 471 621
rect 477 615 483 621
rect 489 615 495 621
rect 501 615 507 621
rect 513 615 519 621
rect 525 615 531 621
rect 537 615 543 621
rect 549 615 555 621
rect 561 615 567 621
rect 573 615 579 621
rect 585 615 591 621
rect 597 615 603 621
rect 609 615 615 621
rect 621 615 627 621
rect 633 615 639 621
rect 645 615 651 621
rect 657 615 663 621
rect 669 615 675 621
rect 681 615 687 621
rect 693 615 699 621
rect 705 615 711 621
rect 717 615 723 621
rect 729 615 735 621
rect 741 615 747 621
rect 753 615 759 621
rect 765 615 771 621
rect 777 615 783 621
rect 789 615 795 621
rect 801 615 807 621
rect 813 615 819 621
rect 825 615 831 621
rect 837 615 843 621
rect 849 615 855 621
rect 861 615 867 621
rect 873 615 879 621
rect 885 615 891 621
rect 897 615 903 621
rect 909 615 915 621
rect 921 615 927 621
rect 933 615 939 621
rect 945 615 951 621
rect 957 615 963 621
rect 969 615 975 621
rect 981 615 987 621
rect 993 615 999 621
rect 1005 615 1011 621
rect 1017 615 1023 621
rect 1029 615 1035 621
rect 1041 615 1047 621
rect 1053 615 1059 621
rect 1065 615 1071 621
rect 1077 615 1083 621
rect 1089 615 1095 621
rect 1101 615 1107 621
rect 1113 615 1119 621
rect 1125 615 1131 621
rect 1137 615 1143 621
rect 1149 615 1155 621
rect 1161 615 1167 621
rect 1173 615 1179 621
rect 1185 615 1191 621
rect 1197 615 1203 621
rect 1209 615 1215 621
rect 1221 615 1227 621
rect 1233 615 1239 621
rect 1245 615 1251 621
rect 1257 615 1263 621
rect 1269 615 1275 621
rect 1281 615 1287 621
rect 1293 615 1299 621
rect 1305 615 1311 621
rect 1317 615 1323 621
rect 1329 615 1335 621
rect 1341 615 1347 621
rect 1353 615 1359 621
rect 1365 615 1371 621
rect 1377 615 1383 621
rect 1389 615 1395 621
rect 1401 615 1407 621
rect 1413 615 1419 621
rect 1425 615 1431 621
rect 1437 615 1443 621
rect 1449 615 1455 621
rect 1461 615 1467 621
rect 1473 615 1479 621
rect 1485 615 1491 621
rect 1497 615 1503 621
rect 1509 615 1515 621
rect 1521 615 1527 621
rect 1533 615 1539 621
rect 1545 615 1551 621
rect 1557 615 1563 621
rect 1569 615 1575 621
rect 1581 615 1587 621
rect 1593 615 1599 621
rect 1605 615 1611 621
rect 1617 615 1623 621
rect 1629 615 1632 621
rect -108 612 1632 615
rect -108 609 -96 612
rect -108 603 -105 609
rect -99 603 -96 609
rect -108 597 -96 603
rect 1620 609 1632 612
rect 1620 603 1623 609
rect 1629 603 1632 609
rect -108 591 -105 597
rect -99 591 -96 597
rect -108 585 -96 591
rect -108 579 -105 585
rect -99 579 -96 585
rect -108 573 -96 579
rect -108 567 -105 573
rect -99 567 -96 573
rect -108 561 -96 567
rect -108 555 -105 561
rect -99 555 -96 561
rect -108 549 -96 555
rect -108 543 -105 549
rect -99 543 -96 549
rect -108 537 -96 543
rect -108 531 -105 537
rect -99 531 -96 537
rect -108 525 -96 531
rect -108 519 -105 525
rect -99 519 -96 525
rect -108 513 -96 519
rect -108 507 -105 513
rect -99 507 -96 513
rect -108 501 -96 507
rect -108 495 -105 501
rect -99 495 -96 501
rect -108 489 -96 495
rect 1620 597 1632 603
rect 1620 591 1623 597
rect 1629 591 1632 597
rect 1620 585 1632 591
rect 1620 579 1623 585
rect 1629 579 1632 585
rect 1620 573 1632 579
rect 1620 567 1623 573
rect 1629 567 1632 573
rect 1620 561 1632 567
rect 1620 555 1623 561
rect 1629 555 1632 561
rect 1620 549 1632 555
rect 1620 543 1623 549
rect 1629 543 1632 549
rect 1620 537 1632 543
rect 1620 531 1623 537
rect 1629 531 1632 537
rect 1620 525 1632 531
rect 1620 519 1623 525
rect 1629 519 1632 525
rect 1620 513 1632 519
rect 1620 507 1623 513
rect 1629 507 1632 513
rect 1620 501 1632 507
rect 1620 495 1623 501
rect 1629 495 1632 501
rect -108 483 -105 489
rect -99 483 -96 489
rect -108 480 -96 483
rect 1620 489 1632 495
rect 1620 483 1623 489
rect 1629 483 1632 489
rect 1620 480 1632 483
rect -108 477 1632 480
rect -108 471 -105 477
rect -99 471 -93 477
rect -87 471 -81 477
rect -75 471 -69 477
rect -63 471 -57 477
rect -51 471 -45 477
rect -39 471 -33 477
rect -27 471 -21 477
rect -15 471 -9 477
rect -3 471 3 477
rect 9 471 15 477
rect 21 471 27 477
rect 33 471 39 477
rect 45 471 51 477
rect 57 471 63 477
rect 69 471 75 477
rect 81 471 87 477
rect 93 471 99 477
rect 105 471 111 477
rect 117 471 123 477
rect 129 471 135 477
rect 141 471 147 477
rect 153 471 159 477
rect 165 471 171 477
rect 177 471 183 477
rect 189 471 195 477
rect 201 471 207 477
rect 213 471 219 477
rect 225 471 231 477
rect 237 471 243 477
rect 249 471 255 477
rect 261 471 267 477
rect 273 471 279 477
rect 285 471 291 477
rect 297 471 303 477
rect 309 471 315 477
rect 321 471 327 477
rect 333 471 339 477
rect 345 471 351 477
rect 357 471 363 477
rect 369 471 375 477
rect 381 471 387 477
rect 393 471 399 477
rect 405 471 411 477
rect 417 471 423 477
rect 429 471 435 477
rect 441 471 447 477
rect 453 471 459 477
rect 465 471 471 477
rect 477 471 483 477
rect 489 471 495 477
rect 501 471 507 477
rect 513 471 519 477
rect 525 471 531 477
rect 537 471 543 477
rect 549 471 555 477
rect 561 471 567 477
rect 573 471 579 477
rect 585 471 591 477
rect 597 471 603 477
rect 609 471 615 477
rect 621 471 627 477
rect 633 471 639 477
rect 645 471 651 477
rect 657 471 663 477
rect 669 471 675 477
rect 681 471 687 477
rect 693 471 699 477
rect 705 471 711 477
rect 717 471 723 477
rect 729 471 735 477
rect 741 471 747 477
rect 753 471 759 477
rect 765 471 771 477
rect 777 471 783 477
rect 789 471 795 477
rect 801 471 807 477
rect 813 471 819 477
rect 825 471 831 477
rect 837 471 843 477
rect 849 471 855 477
rect 861 471 867 477
rect 873 471 879 477
rect 885 471 891 477
rect 897 471 903 477
rect 909 471 915 477
rect 921 471 927 477
rect 933 471 939 477
rect 945 471 951 477
rect 957 471 963 477
rect 969 471 975 477
rect 981 471 987 477
rect 993 471 999 477
rect 1005 471 1011 477
rect 1017 471 1023 477
rect 1029 471 1035 477
rect 1041 471 1047 477
rect 1053 471 1059 477
rect 1065 471 1071 477
rect 1077 471 1083 477
rect 1089 471 1095 477
rect 1101 471 1107 477
rect 1113 471 1119 477
rect 1125 471 1131 477
rect 1137 471 1143 477
rect 1149 471 1155 477
rect 1161 471 1167 477
rect 1173 471 1179 477
rect 1185 471 1191 477
rect 1197 471 1203 477
rect 1209 471 1215 477
rect 1221 471 1227 477
rect 1233 471 1239 477
rect 1245 471 1251 477
rect 1257 471 1263 477
rect 1269 471 1275 477
rect 1281 471 1287 477
rect 1293 471 1299 477
rect 1305 471 1311 477
rect 1317 471 1323 477
rect 1329 471 1335 477
rect 1341 471 1347 477
rect 1353 471 1359 477
rect 1365 471 1371 477
rect 1377 471 1383 477
rect 1389 471 1395 477
rect 1401 471 1407 477
rect 1413 471 1419 477
rect 1425 471 1431 477
rect 1437 471 1443 477
rect 1449 471 1455 477
rect 1461 471 1467 477
rect 1473 471 1479 477
rect 1485 471 1491 477
rect 1497 471 1503 477
rect 1509 471 1515 477
rect 1521 471 1527 477
rect 1533 471 1539 477
rect 1545 471 1551 477
rect 1557 471 1563 477
rect 1569 471 1575 477
rect 1581 471 1587 477
rect 1593 471 1599 477
rect 1605 471 1611 477
rect 1617 471 1623 477
rect 1629 471 1632 477
rect -108 468 1632 471
rect -108 465 -96 468
rect -108 459 -105 465
rect -99 459 -96 465
rect -108 453 -96 459
rect 1620 465 1632 468
rect 1620 459 1623 465
rect 1629 459 1632 465
rect -108 447 -105 453
rect -99 447 -96 453
rect -108 441 -96 447
rect -108 435 -105 441
rect -99 435 -96 441
rect -108 429 -96 435
rect -108 423 -105 429
rect -99 423 -96 429
rect -108 417 -96 423
rect -108 411 -105 417
rect -99 411 -96 417
rect -108 405 -96 411
rect -108 399 -105 405
rect -99 399 -96 405
rect -108 393 -96 399
rect -108 387 -105 393
rect -99 387 -96 393
rect -108 381 -96 387
rect -108 375 -105 381
rect -99 375 -96 381
rect -108 369 -96 375
rect -108 363 -105 369
rect -99 363 -96 369
rect -108 357 -96 363
rect -108 351 -105 357
rect -99 351 -96 357
rect -108 345 -96 351
rect 1620 453 1632 459
rect 1620 447 1623 453
rect 1629 447 1632 453
rect 1620 441 1632 447
rect 1620 435 1623 441
rect 1629 435 1632 441
rect 1620 429 1632 435
rect 1620 423 1623 429
rect 1629 423 1632 429
rect 1620 417 1632 423
rect 1620 411 1623 417
rect 1629 411 1632 417
rect 1620 405 1632 411
rect 1620 399 1623 405
rect 1629 399 1632 405
rect 1620 393 1632 399
rect 1620 387 1623 393
rect 1629 387 1632 393
rect 1620 381 1632 387
rect 1620 375 1623 381
rect 1629 375 1632 381
rect 1620 369 1632 375
rect 1620 363 1623 369
rect 1629 363 1632 369
rect 1620 357 1632 363
rect 1620 351 1623 357
rect 1629 351 1632 357
rect -108 339 -105 345
rect -99 339 -96 345
rect -108 336 -96 339
rect 1620 345 1632 351
rect 1620 339 1623 345
rect 1629 339 1632 345
rect 1620 336 1632 339
rect -108 333 1632 336
rect -108 327 -105 333
rect -99 327 -93 333
rect -87 327 -81 333
rect -75 327 -69 333
rect -63 327 -57 333
rect -51 327 -45 333
rect -39 327 -33 333
rect -27 327 -21 333
rect -15 327 -9 333
rect -3 327 3 333
rect 9 327 15 333
rect 21 327 27 333
rect 33 327 39 333
rect 45 327 51 333
rect 57 327 63 333
rect 69 327 75 333
rect 81 327 87 333
rect 93 327 99 333
rect 105 327 111 333
rect 117 327 123 333
rect 129 327 135 333
rect 141 327 147 333
rect 153 327 159 333
rect 165 327 171 333
rect 177 327 183 333
rect 189 327 195 333
rect 201 327 207 333
rect 213 327 219 333
rect 225 327 231 333
rect 237 327 243 333
rect 249 327 255 333
rect 261 327 267 333
rect 273 327 279 333
rect 285 327 291 333
rect 297 327 303 333
rect 309 327 315 333
rect 321 327 327 333
rect 333 327 339 333
rect 345 327 351 333
rect 357 327 363 333
rect 369 327 375 333
rect 381 327 387 333
rect 393 327 399 333
rect 405 327 411 333
rect 417 327 423 333
rect 429 327 435 333
rect 441 327 447 333
rect 453 327 459 333
rect 465 327 471 333
rect 477 327 483 333
rect 489 327 495 333
rect 501 327 507 333
rect 513 327 519 333
rect 525 327 531 333
rect 537 327 543 333
rect 549 327 555 333
rect 561 327 567 333
rect 573 327 579 333
rect 585 327 591 333
rect 597 327 603 333
rect 609 327 615 333
rect 621 327 627 333
rect 633 327 639 333
rect 645 327 651 333
rect 657 327 663 333
rect 669 327 675 333
rect 681 327 687 333
rect 693 327 699 333
rect 705 327 711 333
rect 717 327 723 333
rect 729 327 735 333
rect 741 327 747 333
rect 753 327 759 333
rect 765 327 771 333
rect 777 327 783 333
rect 789 327 795 333
rect 801 327 807 333
rect 813 327 819 333
rect 825 327 831 333
rect 837 327 843 333
rect 849 327 855 333
rect 861 327 867 333
rect 873 327 879 333
rect 885 327 891 333
rect 897 327 903 333
rect 909 327 915 333
rect 921 327 927 333
rect 933 327 939 333
rect 945 327 951 333
rect 957 327 963 333
rect 969 327 975 333
rect 981 327 987 333
rect 993 327 999 333
rect 1005 327 1011 333
rect 1017 327 1023 333
rect 1029 327 1035 333
rect 1041 327 1047 333
rect 1053 327 1059 333
rect 1065 327 1071 333
rect 1077 327 1083 333
rect 1089 327 1095 333
rect 1101 327 1107 333
rect 1113 327 1119 333
rect 1125 327 1131 333
rect 1137 327 1143 333
rect 1149 327 1155 333
rect 1161 327 1167 333
rect 1173 327 1179 333
rect 1185 327 1191 333
rect 1197 327 1203 333
rect 1209 327 1215 333
rect 1221 327 1227 333
rect 1233 327 1239 333
rect 1245 327 1251 333
rect 1257 327 1263 333
rect 1269 327 1275 333
rect 1281 327 1287 333
rect 1293 327 1299 333
rect 1305 327 1311 333
rect 1317 327 1323 333
rect 1329 327 1335 333
rect 1341 327 1347 333
rect 1353 327 1359 333
rect 1365 327 1371 333
rect 1377 327 1383 333
rect 1389 327 1395 333
rect 1401 327 1407 333
rect 1413 327 1419 333
rect 1425 327 1431 333
rect 1437 327 1443 333
rect 1449 327 1455 333
rect 1461 327 1467 333
rect 1473 327 1479 333
rect 1485 327 1491 333
rect 1497 327 1503 333
rect 1509 327 1515 333
rect 1521 327 1527 333
rect 1533 327 1539 333
rect 1545 327 1551 333
rect 1557 327 1563 333
rect 1569 327 1575 333
rect 1581 327 1587 333
rect 1593 327 1599 333
rect 1605 327 1611 333
rect 1617 327 1623 333
rect 1629 327 1632 333
rect -108 324 1632 327
rect -108 321 -96 324
rect -108 315 -105 321
rect -99 315 -96 321
rect -108 309 -96 315
rect -108 303 -105 309
rect -99 303 -96 309
rect -108 297 -96 303
rect -108 291 -105 297
rect -99 291 -96 297
rect -108 285 -96 291
rect -108 279 -105 285
rect -99 279 -96 285
rect -108 273 -96 279
rect -108 267 -105 273
rect -99 267 -96 273
rect -108 261 -96 267
rect -108 255 -105 261
rect -99 255 -96 261
rect -108 249 -96 255
rect -108 243 -105 249
rect -99 243 -96 249
rect -108 237 -96 243
rect -108 231 -105 237
rect -99 231 -96 237
rect -108 225 -96 231
rect -108 219 -105 225
rect -99 219 -96 225
rect -108 213 -96 219
rect -108 207 -105 213
rect -99 207 -96 213
rect -108 201 -96 207
rect -108 195 -105 201
rect -99 195 -96 201
rect -108 189 -96 195
rect -108 183 -105 189
rect -99 183 -96 189
rect -108 177 -96 183
rect -108 171 -105 177
rect -99 171 -96 177
rect -108 165 -96 171
rect -108 159 -105 165
rect -99 159 -96 165
rect -108 153 -96 159
rect -108 147 -105 153
rect -99 147 -96 153
rect -108 141 -96 147
rect -108 135 -105 141
rect -99 135 -96 141
rect -108 129 -96 135
rect -108 123 -105 129
rect -99 123 -96 129
rect -108 117 -96 123
rect -108 111 -105 117
rect -99 111 -96 117
rect -108 105 -96 111
rect -108 99 -105 105
rect -99 99 -96 105
rect -108 96 -96 99
rect 1620 321 1632 324
rect 1620 315 1623 321
rect 1629 315 1632 321
rect 1620 309 1632 315
rect 1620 303 1623 309
rect 1629 303 1632 309
rect 1620 297 1632 303
rect 1620 291 1623 297
rect 1629 291 1632 297
rect 1620 285 1632 291
rect 1620 279 1623 285
rect 1629 279 1632 285
rect 1620 273 1632 279
rect 1620 267 1623 273
rect 1629 267 1632 273
rect 1620 261 1632 267
rect 1620 255 1623 261
rect 1629 255 1632 261
rect 1620 249 1632 255
rect 1620 243 1623 249
rect 1629 243 1632 249
rect 1620 237 1632 243
rect 1620 231 1623 237
rect 1629 231 1632 237
rect 1620 225 1632 231
rect 1620 219 1623 225
rect 1629 219 1632 225
rect 1620 213 1632 219
rect 1620 207 1623 213
rect 1629 207 1632 213
rect 1620 201 1632 207
rect 1620 195 1623 201
rect 1629 195 1632 201
rect 1620 189 1632 195
rect 1620 183 1623 189
rect 1629 183 1632 189
rect 1620 177 1632 183
rect 1620 171 1623 177
rect 1629 171 1632 177
rect 1620 165 1632 171
rect 1620 159 1623 165
rect 1629 159 1632 165
rect 1620 153 1632 159
rect 1620 147 1623 153
rect 1629 147 1632 153
rect 1620 141 1632 147
rect 1620 135 1623 141
rect 1629 135 1632 141
rect 1620 129 1632 135
rect 1620 123 1623 129
rect 1629 123 1632 129
rect 1620 117 1632 123
rect 1620 111 1623 117
rect 1629 111 1632 117
rect 1620 105 1632 111
rect 1620 99 1623 105
rect 1629 99 1632 105
rect 1620 96 1632 99
rect -108 93 1632 96
rect -108 87 -105 93
rect -99 87 -93 93
rect -87 87 -81 93
rect -75 87 -69 93
rect -63 87 -57 93
rect -51 87 -45 93
rect -39 87 -33 93
rect -27 87 -21 93
rect -15 87 -9 93
rect -3 87 3 93
rect 9 87 15 93
rect 21 87 27 93
rect 33 87 39 93
rect 45 87 51 93
rect 57 87 63 93
rect 69 87 75 93
rect 81 87 87 93
rect 93 87 99 93
rect 105 87 111 93
rect 117 87 123 93
rect 129 87 135 93
rect 141 87 147 93
rect 153 87 159 93
rect 165 87 171 93
rect 177 87 183 93
rect 189 87 195 93
rect 201 87 207 93
rect 213 87 219 93
rect 225 87 231 93
rect 237 87 243 93
rect 249 87 255 93
rect 261 87 267 93
rect 273 87 279 93
rect 285 87 291 93
rect 297 87 303 93
rect 309 87 315 93
rect 321 87 327 93
rect 333 87 339 93
rect 345 87 351 93
rect 357 87 363 93
rect 369 87 375 93
rect 381 87 387 93
rect 393 87 399 93
rect 405 87 411 93
rect 417 87 423 93
rect 429 87 435 93
rect 441 87 447 93
rect 453 87 459 93
rect 465 87 471 93
rect 477 87 483 93
rect 489 87 495 93
rect 501 87 507 93
rect 513 87 519 93
rect 525 87 531 93
rect 537 87 543 93
rect 549 87 555 93
rect 561 87 567 93
rect 573 87 579 93
rect 585 87 591 93
rect 597 87 603 93
rect 609 87 615 93
rect 621 87 627 93
rect 633 87 639 93
rect 645 87 651 93
rect 657 87 663 93
rect 669 87 675 93
rect 681 87 687 93
rect 693 87 699 93
rect 705 87 711 93
rect 717 87 723 93
rect 729 87 735 93
rect 741 87 747 93
rect 753 87 759 93
rect 765 87 771 93
rect 777 87 783 93
rect 789 87 795 93
rect 801 87 807 93
rect 813 87 819 93
rect 825 87 831 93
rect 837 87 843 93
rect 849 87 855 93
rect 861 87 867 93
rect 873 87 879 93
rect 885 87 891 93
rect 897 87 903 93
rect 909 87 915 93
rect 921 87 927 93
rect 933 87 939 93
rect 945 87 951 93
rect 957 87 963 93
rect 969 87 975 93
rect 981 87 987 93
rect 993 87 999 93
rect 1005 87 1011 93
rect 1017 87 1023 93
rect 1029 87 1035 93
rect 1041 87 1047 93
rect 1053 87 1059 93
rect 1065 87 1071 93
rect 1077 87 1083 93
rect 1089 87 1095 93
rect 1101 87 1107 93
rect 1113 87 1119 93
rect 1125 87 1131 93
rect 1137 87 1143 93
rect 1149 87 1155 93
rect 1161 87 1167 93
rect 1173 87 1179 93
rect 1185 87 1191 93
rect 1197 87 1203 93
rect 1209 87 1215 93
rect 1221 87 1227 93
rect 1233 87 1239 93
rect 1245 87 1251 93
rect 1257 87 1263 93
rect 1269 87 1275 93
rect 1281 87 1287 93
rect 1293 87 1299 93
rect 1305 87 1311 93
rect 1317 87 1323 93
rect 1329 87 1335 93
rect 1341 87 1347 93
rect 1353 87 1359 93
rect 1365 87 1371 93
rect 1377 87 1383 93
rect 1389 87 1395 93
rect 1401 87 1407 93
rect 1413 87 1419 93
rect 1425 87 1431 93
rect 1437 87 1443 93
rect 1449 87 1455 93
rect 1461 87 1467 93
rect 1473 87 1479 93
rect 1485 87 1491 93
rect 1497 87 1503 93
rect 1509 87 1515 93
rect 1521 87 1527 93
rect 1533 87 1539 93
rect 1545 87 1551 93
rect 1557 87 1563 93
rect 1569 87 1575 93
rect 1581 87 1587 93
rect 1593 87 1599 93
rect 1605 87 1611 93
rect 1617 87 1623 93
rect 1629 87 1632 93
rect -108 84 1632 87
rect -108 81 -96 84
rect -108 75 -105 81
rect -99 75 -96 81
rect -108 69 -96 75
rect 1620 81 1632 84
rect 1620 75 1623 81
rect 1629 75 1632 81
rect -108 63 -105 69
rect -99 63 -96 69
rect -108 57 -96 63
rect -108 51 -105 57
rect -99 51 -96 57
rect -108 45 -96 51
rect 1620 69 1632 75
rect 1620 63 1623 69
rect 1629 63 1632 69
rect 1620 57 1632 63
rect 1620 51 1623 57
rect 1629 51 1632 57
rect -108 39 -105 45
rect -99 39 -96 45
rect -108 33 -96 39
rect -108 27 -105 33
rect -99 27 -96 33
rect -108 21 -96 27
rect -108 15 -105 21
rect -99 15 -96 21
rect -108 9 -96 15
rect 1620 45 1632 51
rect 1620 39 1623 45
rect 1629 39 1632 45
rect 1620 33 1632 39
rect 1620 27 1623 33
rect 1629 27 1632 33
rect 1620 21 1632 27
rect 1620 15 1623 21
rect 1629 15 1632 21
rect -108 3 -105 9
rect -99 3 -96 9
rect 1620 9 1632 15
rect -108 0 -96 3
rect 1620 3 1623 9
rect 1629 3 1632 9
rect 1620 0 1632 3
rect -108 -3 1632 0
rect -108 -9 -105 -3
rect -99 -9 -93 -3
rect -87 -9 -81 -3
rect -75 -9 -69 -3
rect -63 -9 -57 -3
rect -51 -9 -45 -3
rect -39 -9 -33 -3
rect -27 -9 -21 -3
rect -15 -9 -9 -3
rect -3 -9 3 -3
rect 9 -9 15 -3
rect 21 -9 27 -3
rect 33 -9 39 -3
rect 45 -9 51 -3
rect 57 -9 63 -3
rect 69 -9 75 -3
rect 81 -9 87 -3
rect 93 -9 99 -3
rect 105 -9 111 -3
rect 117 -9 123 -3
rect 129 -9 135 -3
rect 141 -9 147 -3
rect 153 -9 159 -3
rect 165 -9 171 -3
rect 177 -9 183 -3
rect 189 -9 195 -3
rect 201 -9 207 -3
rect 213 -9 219 -3
rect 225 -9 231 -3
rect 237 -9 243 -3
rect 249 -9 255 -3
rect 261 -9 267 -3
rect 273 -9 279 -3
rect 285 -9 291 -3
rect 297 -9 303 -3
rect 309 -9 315 -3
rect 321 -9 327 -3
rect 333 -9 339 -3
rect 345 -9 351 -3
rect 357 -9 363 -3
rect 369 -9 375 -3
rect 381 -9 387 -3
rect 393 -9 399 -3
rect 405 -9 411 -3
rect 417 -9 423 -3
rect 429 -9 435 -3
rect 441 -9 447 -3
rect 453 -9 459 -3
rect 465 -9 471 -3
rect 477 -9 483 -3
rect 489 -9 495 -3
rect 501 -9 507 -3
rect 513 -9 519 -3
rect 525 -9 531 -3
rect 537 -9 543 -3
rect 549 -9 555 -3
rect 561 -9 567 -3
rect 573 -9 579 -3
rect 585 -9 591 -3
rect 597 -9 603 -3
rect 609 -9 615 -3
rect 621 -9 627 -3
rect 633 -9 639 -3
rect 645 -9 651 -3
rect 657 -9 663 -3
rect 669 -9 675 -3
rect 681 -9 687 -3
rect 693 -9 699 -3
rect 705 -9 711 -3
rect 717 -9 723 -3
rect 729 -9 735 -3
rect 741 -9 747 -3
rect 753 -9 759 -3
rect 765 -9 771 -3
rect 777 -9 783 -3
rect 789 -9 795 -3
rect 801 -9 807 -3
rect 813 -9 819 -3
rect 825 -9 831 -3
rect 837 -9 843 -3
rect 849 -9 855 -3
rect 861 -9 867 -3
rect 873 -9 879 -3
rect 885 -9 891 -3
rect 897 -9 903 -3
rect 909 -9 915 -3
rect 921 -9 927 -3
rect 933 -9 939 -3
rect 945 -9 951 -3
rect 957 -9 963 -3
rect 969 -9 975 -3
rect 981 -9 987 -3
rect 993 -9 999 -3
rect 1005 -9 1011 -3
rect 1017 -9 1023 -3
rect 1029 -9 1035 -3
rect 1041 -9 1047 -3
rect 1053 -9 1059 -3
rect 1065 -9 1071 -3
rect 1077 -9 1083 -3
rect 1089 -9 1095 -3
rect 1101 -9 1107 -3
rect 1113 -9 1119 -3
rect 1125 -9 1131 -3
rect 1137 -9 1143 -3
rect 1149 -9 1155 -3
rect 1161 -9 1167 -3
rect 1173 -9 1179 -3
rect 1185 -9 1191 -3
rect 1197 -9 1203 -3
rect 1209 -9 1215 -3
rect 1221 -9 1227 -3
rect 1233 -9 1239 -3
rect 1245 -9 1251 -3
rect 1257 -9 1263 -3
rect 1269 -9 1275 -3
rect 1281 -9 1287 -3
rect 1293 -9 1299 -3
rect 1305 -9 1311 -3
rect 1317 -9 1323 -3
rect 1329 -9 1335 -3
rect 1341 -9 1347 -3
rect 1353 -9 1359 -3
rect 1365 -9 1371 -3
rect 1377 -9 1383 -3
rect 1389 -9 1395 -3
rect 1401 -9 1407 -3
rect 1413 -9 1419 -3
rect 1425 -9 1431 -3
rect 1437 -9 1443 -3
rect 1449 -9 1455 -3
rect 1461 -9 1467 -3
rect 1473 -9 1479 -3
rect 1485 -9 1491 -3
rect 1497 -9 1503 -3
rect 1509 -9 1515 -3
rect 1521 -9 1527 -3
rect 1533 -9 1539 -3
rect 1545 -9 1551 -3
rect 1557 -9 1563 -3
rect 1569 -9 1575 -3
rect 1581 -9 1587 -3
rect 1593 -9 1599 -3
rect 1605 -9 1611 -3
rect 1617 -9 1623 -3
rect 1629 -9 1632 -3
rect -108 -12 1632 -9
rect -108 -15 -96 -12
rect -108 -21 -105 -15
rect -99 -21 -96 -15
rect -108 -27 -96 -21
rect -108 -33 -105 -27
rect -99 -33 -96 -27
rect -108 -39 -96 -33
rect -108 -45 -105 -39
rect -99 -45 -96 -39
rect -108 -51 -96 -45
rect -108 -57 -105 -51
rect -99 -57 -96 -51
rect -108 -63 -96 -57
rect -108 -69 -105 -63
rect -99 -69 -96 -63
rect -108 -75 -96 -69
rect -108 -81 -105 -75
rect -99 -81 -96 -75
rect -108 -87 -96 -81
rect -108 -93 -105 -87
rect -99 -93 -96 -87
rect -108 -99 -96 -93
rect -108 -105 -105 -99
rect -99 -105 -96 -99
rect -108 -111 -96 -105
rect -108 -117 -105 -111
rect -99 -117 -96 -111
rect -108 -123 -96 -117
rect -108 -129 -105 -123
rect -99 -129 -96 -123
rect -108 -135 -96 -129
rect -108 -141 -105 -135
rect -99 -141 -96 -135
rect -108 -147 -96 -141
rect -108 -153 -105 -147
rect -99 -153 -96 -147
rect -108 -159 -96 -153
rect -108 -165 -105 -159
rect -99 -165 -96 -159
rect -108 -171 -96 -165
rect -108 -177 -105 -171
rect -99 -177 -96 -171
rect -108 -183 -96 -177
rect -108 -189 -105 -183
rect -99 -189 -96 -183
rect -108 -192 -96 -189
rect 1620 -15 1632 -12
rect 1620 -21 1623 -15
rect 1629 -21 1632 -15
rect 1620 -27 1632 -21
rect 1620 -33 1623 -27
rect 1629 -33 1632 -27
rect 1620 -39 1632 -33
rect 1620 -45 1623 -39
rect 1629 -45 1632 -39
rect 1620 -51 1632 -45
rect 1620 -57 1623 -51
rect 1629 -57 1632 -51
rect 1620 -63 1632 -57
rect 1620 -69 1623 -63
rect 1629 -69 1632 -63
rect 1620 -75 1632 -69
rect 1620 -81 1623 -75
rect 1629 -81 1632 -75
rect 1620 -87 1632 -81
rect 1620 -93 1623 -87
rect 1629 -93 1632 -87
rect 1620 -99 1632 -93
rect 1620 -105 1623 -99
rect 1629 -105 1632 -99
rect 1620 -111 1632 -105
rect 1620 -117 1623 -111
rect 1629 -117 1632 -111
rect 1620 -123 1632 -117
rect 1620 -129 1623 -123
rect 1629 -129 1632 -123
rect 1620 -135 1632 -129
rect 1620 -141 1623 -135
rect 1629 -141 1632 -135
rect 1620 -147 1632 -141
rect 1620 -153 1623 -147
rect 1629 -153 1632 -147
rect 1620 -159 1632 -153
rect 1620 -165 1623 -159
rect 1629 -165 1632 -159
rect 1620 -171 1632 -165
rect 1620 -177 1623 -171
rect 1629 -177 1632 -171
rect 1620 -183 1632 -177
rect 1620 -189 1623 -183
rect 1629 -189 1632 -183
rect 1620 -192 1632 -189
rect -108 -195 1632 -192
rect -108 -201 -105 -195
rect -99 -201 -93 -195
rect -87 -201 -81 -195
rect -75 -201 -69 -195
rect -63 -201 -57 -195
rect -51 -201 -45 -195
rect -39 -201 -33 -195
rect -27 -201 -21 -195
rect -15 -201 -9 -195
rect -3 -201 3 -195
rect 9 -201 15 -195
rect 21 -201 27 -195
rect 33 -201 39 -195
rect 45 -201 51 -195
rect 57 -201 63 -195
rect 69 -201 75 -195
rect 81 -201 87 -195
rect 93 -201 99 -195
rect 105 -201 111 -195
rect 117 -201 123 -195
rect 129 -201 135 -195
rect 141 -201 147 -195
rect 153 -201 159 -195
rect 165 -201 171 -195
rect 177 -201 183 -195
rect 189 -201 195 -195
rect 201 -201 207 -195
rect 213 -201 219 -195
rect 225 -201 231 -195
rect 237 -201 243 -195
rect 249 -201 255 -195
rect 261 -201 267 -195
rect 273 -201 279 -195
rect 285 -201 291 -195
rect 297 -201 303 -195
rect 309 -201 315 -195
rect 321 -201 327 -195
rect 333 -201 339 -195
rect 345 -201 351 -195
rect 357 -201 363 -195
rect 369 -201 375 -195
rect 381 -201 387 -195
rect 393 -201 399 -195
rect 405 -201 411 -195
rect 417 -201 423 -195
rect 429 -201 435 -195
rect 441 -201 447 -195
rect 453 -201 459 -195
rect 465 -201 471 -195
rect 477 -201 483 -195
rect 489 -201 495 -195
rect 501 -201 507 -195
rect 513 -201 519 -195
rect 525 -201 531 -195
rect 537 -201 543 -195
rect 549 -201 555 -195
rect 561 -201 567 -195
rect 573 -201 579 -195
rect 585 -201 591 -195
rect 597 -201 603 -195
rect 609 -201 615 -195
rect 621 -201 627 -195
rect 633 -201 639 -195
rect 645 -201 651 -195
rect 657 -201 663 -195
rect 669 -201 675 -195
rect 681 -201 687 -195
rect 693 -201 699 -195
rect 705 -201 711 -195
rect 717 -201 723 -195
rect 729 -201 735 -195
rect 741 -201 747 -195
rect 753 -201 759 -195
rect 765 -201 771 -195
rect 777 -201 783 -195
rect 789 -201 795 -195
rect 801 -201 807 -195
rect 813 -201 819 -195
rect 825 -201 831 -195
rect 837 -201 843 -195
rect 849 -201 855 -195
rect 861 -201 867 -195
rect 873 -201 879 -195
rect 885 -201 891 -195
rect 897 -201 903 -195
rect 909 -201 915 -195
rect 921 -201 927 -195
rect 933 -201 939 -195
rect 945 -201 951 -195
rect 957 -201 963 -195
rect 969 -201 975 -195
rect 981 -201 987 -195
rect 993 -201 999 -195
rect 1005 -201 1011 -195
rect 1017 -201 1023 -195
rect 1029 -201 1035 -195
rect 1041 -201 1047 -195
rect 1053 -201 1059 -195
rect 1065 -201 1071 -195
rect 1077 -201 1083 -195
rect 1089 -201 1095 -195
rect 1101 -201 1107 -195
rect 1113 -201 1119 -195
rect 1125 -201 1131 -195
rect 1137 -201 1143 -195
rect 1149 -201 1155 -195
rect 1161 -201 1167 -195
rect 1173 -201 1179 -195
rect 1185 -201 1191 -195
rect 1197 -201 1203 -195
rect 1209 -201 1215 -195
rect 1221 -201 1227 -195
rect 1233 -201 1239 -195
rect 1245 -201 1251 -195
rect 1257 -201 1263 -195
rect 1269 -201 1275 -195
rect 1281 -201 1287 -195
rect 1293 -201 1299 -195
rect 1305 -201 1311 -195
rect 1317 -201 1323 -195
rect 1329 -201 1335 -195
rect 1341 -201 1347 -195
rect 1353 -201 1359 -195
rect 1365 -201 1371 -195
rect 1377 -201 1383 -195
rect 1389 -201 1395 -195
rect 1401 -201 1407 -195
rect 1413 -201 1419 -195
rect 1425 -201 1431 -195
rect 1437 -201 1443 -195
rect 1449 -201 1455 -195
rect 1461 -201 1563 -195
rect 1569 -201 1575 -195
rect 1581 -201 1587 -195
rect 1593 -201 1599 -195
rect 1605 -201 1611 -195
rect 1617 -201 1623 -195
rect 1629 -201 1632 -195
rect -108 -204 1632 -201
<< nsubdiff >>
rect -84 597 1608 600
rect -84 591 -81 597
rect -75 591 -69 597
rect -63 591 -57 597
rect -51 591 -45 597
rect -39 591 -33 597
rect -27 591 -21 597
rect -15 591 -9 597
rect -3 591 3 597
rect 9 591 15 597
rect 21 591 27 597
rect 33 591 39 597
rect 45 591 51 597
rect 57 591 63 597
rect 69 591 75 597
rect 81 591 87 597
rect 93 591 99 597
rect 105 591 111 597
rect 117 591 123 597
rect 129 591 135 597
rect 141 591 147 597
rect 153 591 159 597
rect 165 591 171 597
rect 177 591 183 597
rect 189 591 195 597
rect 201 591 207 597
rect 213 591 219 597
rect 225 591 231 597
rect 237 591 243 597
rect 249 591 255 597
rect 261 591 267 597
rect 273 591 279 597
rect 285 591 291 597
rect 297 591 303 597
rect 309 591 315 597
rect 321 591 327 597
rect 333 591 339 597
rect 345 591 351 597
rect 357 591 363 597
rect 369 591 375 597
rect 381 591 387 597
rect 393 591 399 597
rect 405 591 411 597
rect 417 591 423 597
rect 429 591 435 597
rect 441 591 447 597
rect 453 591 459 597
rect 465 591 471 597
rect 477 591 483 597
rect 489 591 495 597
rect 501 591 507 597
rect 513 591 519 597
rect 525 591 531 597
rect 537 591 543 597
rect 549 591 555 597
rect 561 591 567 597
rect 573 591 579 597
rect 585 591 591 597
rect 597 591 603 597
rect 609 591 615 597
rect 621 591 627 597
rect 633 591 639 597
rect 645 591 651 597
rect 657 591 663 597
rect 669 591 675 597
rect 681 591 687 597
rect 693 591 699 597
rect 705 591 711 597
rect 717 591 723 597
rect 729 591 735 597
rect 741 591 747 597
rect 753 591 759 597
rect 765 591 771 597
rect 777 591 783 597
rect 789 591 795 597
rect 801 591 807 597
rect 813 591 819 597
rect 825 591 831 597
rect 837 591 843 597
rect 849 591 855 597
rect 861 591 867 597
rect 873 591 879 597
rect 885 591 891 597
rect 897 591 903 597
rect 909 591 915 597
rect 921 591 927 597
rect 933 591 939 597
rect 945 591 951 597
rect 957 591 963 597
rect 969 591 975 597
rect 981 591 987 597
rect 993 591 999 597
rect 1005 591 1011 597
rect 1017 591 1023 597
rect 1029 591 1035 597
rect 1041 591 1047 597
rect 1053 591 1059 597
rect 1065 591 1071 597
rect 1077 591 1083 597
rect 1089 591 1095 597
rect 1101 591 1107 597
rect 1113 591 1119 597
rect 1125 591 1131 597
rect 1137 591 1143 597
rect 1149 591 1155 597
rect 1161 591 1167 597
rect 1173 591 1179 597
rect 1185 591 1191 597
rect 1197 591 1203 597
rect 1209 591 1215 597
rect 1221 591 1227 597
rect 1233 591 1239 597
rect 1245 591 1251 597
rect 1257 591 1263 597
rect 1269 591 1275 597
rect 1281 591 1287 597
rect 1293 591 1299 597
rect 1305 591 1311 597
rect 1317 591 1323 597
rect 1329 591 1335 597
rect 1341 591 1347 597
rect 1353 591 1359 597
rect 1365 591 1371 597
rect 1377 591 1383 597
rect 1389 591 1395 597
rect 1401 591 1407 597
rect 1413 591 1419 597
rect 1425 591 1431 597
rect 1437 591 1443 597
rect 1449 591 1455 597
rect 1461 591 1467 597
rect 1473 591 1479 597
rect 1485 591 1491 597
rect 1497 591 1503 597
rect 1509 591 1515 597
rect 1521 591 1527 597
rect 1533 591 1539 597
rect 1545 591 1551 597
rect 1557 591 1563 597
rect 1569 591 1575 597
rect 1581 591 1587 597
rect 1593 591 1599 597
rect 1605 591 1608 597
rect -84 588 1608 591
rect -84 585 -72 588
rect -84 579 -81 585
rect -75 579 -72 585
rect -84 573 -72 579
rect 1596 585 1608 588
rect 1596 579 1599 585
rect 1605 579 1608 585
rect -84 567 -81 573
rect -75 567 -72 573
rect -84 561 -72 567
rect -84 555 -81 561
rect -75 555 -72 561
rect -84 549 -72 555
rect 1596 573 1608 579
rect 1596 567 1599 573
rect 1605 567 1608 573
rect 1596 561 1608 567
rect 1596 555 1599 561
rect 1605 555 1608 561
rect -84 543 -81 549
rect -75 543 -72 549
rect -84 537 -72 543
rect -84 531 -81 537
rect -75 531 -72 537
rect -84 525 -72 531
rect -84 519 -81 525
rect -75 519 -72 525
rect -84 513 -72 519
rect 1596 549 1608 555
rect 1596 543 1599 549
rect 1605 543 1608 549
rect 1596 537 1608 543
rect 1596 531 1599 537
rect 1605 531 1608 537
rect 1596 525 1608 531
rect 1596 519 1599 525
rect 1605 519 1608 525
rect -84 507 -81 513
rect -75 507 -72 513
rect 1596 513 1608 519
rect -84 504 -72 507
rect 1596 507 1599 513
rect 1605 507 1608 513
rect 1596 504 1608 507
rect -84 501 -60 504
rect 1584 501 1608 504
rect -84 495 -81 501
rect -75 495 -69 501
rect -63 495 -60 501
rect 1584 495 1587 501
rect 1593 495 1599 501
rect 1605 495 1608 501
rect -84 492 -60 495
rect 1584 492 1608 495
rect -84 453 1608 456
rect -84 447 -81 453
rect -75 447 -69 453
rect -63 447 -57 453
rect -51 447 -45 453
rect -39 447 -33 453
rect -27 447 -21 453
rect -15 447 -9 453
rect -3 447 3 453
rect 9 447 15 453
rect 21 447 27 453
rect 33 447 39 453
rect 45 447 51 453
rect 57 447 63 453
rect 69 447 75 453
rect 81 447 87 453
rect 93 447 99 453
rect 105 447 111 453
rect 117 447 123 453
rect 129 447 135 453
rect 141 447 147 453
rect 153 447 159 453
rect 165 447 171 453
rect 177 447 183 453
rect 189 447 195 453
rect 201 447 207 453
rect 213 447 219 453
rect 225 447 231 453
rect 237 447 243 453
rect 249 447 255 453
rect 261 447 267 453
rect 273 447 279 453
rect 285 447 291 453
rect 297 447 303 453
rect 309 447 315 453
rect 321 447 327 453
rect 333 447 339 453
rect 345 447 351 453
rect 357 447 363 453
rect 369 447 375 453
rect 381 447 387 453
rect 393 447 399 453
rect 405 447 411 453
rect 417 447 423 453
rect 429 447 435 453
rect 441 447 447 453
rect 453 447 459 453
rect 465 447 471 453
rect 477 447 483 453
rect 489 447 495 453
rect 501 447 507 453
rect 513 447 519 453
rect 525 447 531 453
rect 537 447 543 453
rect 549 447 555 453
rect 561 447 567 453
rect 573 447 579 453
rect 585 447 591 453
rect 597 447 603 453
rect 609 447 615 453
rect 621 447 627 453
rect 633 447 639 453
rect 645 447 651 453
rect 657 447 663 453
rect 669 447 675 453
rect 681 447 687 453
rect 693 447 699 453
rect 705 447 711 453
rect 717 447 723 453
rect 729 447 735 453
rect 741 447 747 453
rect 753 447 759 453
rect 765 447 771 453
rect 777 447 783 453
rect 789 447 795 453
rect 801 447 807 453
rect 813 447 819 453
rect 825 447 831 453
rect 837 447 843 453
rect 849 447 855 453
rect 861 447 867 453
rect 873 447 879 453
rect 885 447 891 453
rect 897 447 903 453
rect 909 447 915 453
rect 921 447 927 453
rect 933 447 939 453
rect 945 447 951 453
rect 957 447 963 453
rect 969 447 975 453
rect 981 447 987 453
rect 993 447 999 453
rect 1005 447 1011 453
rect 1017 447 1023 453
rect 1029 447 1035 453
rect 1041 447 1047 453
rect 1053 447 1059 453
rect 1065 447 1071 453
rect 1077 447 1083 453
rect 1089 447 1095 453
rect 1101 447 1107 453
rect 1113 447 1119 453
rect 1125 447 1131 453
rect 1137 447 1143 453
rect 1149 447 1155 453
rect 1161 447 1167 453
rect 1173 447 1179 453
rect 1185 447 1191 453
rect 1197 447 1203 453
rect 1209 447 1215 453
rect 1221 447 1227 453
rect 1233 447 1239 453
rect 1245 447 1251 453
rect 1257 447 1263 453
rect 1269 447 1275 453
rect 1281 447 1287 453
rect 1293 447 1299 453
rect 1305 447 1311 453
rect 1317 447 1323 453
rect 1329 447 1335 453
rect 1341 447 1347 453
rect 1353 447 1359 453
rect 1365 447 1371 453
rect 1377 447 1383 453
rect 1389 447 1395 453
rect 1401 447 1407 453
rect 1413 447 1419 453
rect 1425 447 1431 453
rect 1437 447 1443 453
rect 1449 447 1455 453
rect 1461 447 1467 453
rect 1473 447 1479 453
rect 1485 447 1491 453
rect 1497 447 1503 453
rect 1509 447 1515 453
rect 1521 447 1527 453
rect 1533 447 1539 453
rect 1545 447 1551 453
rect 1557 447 1563 453
rect 1569 447 1575 453
rect 1581 447 1587 453
rect 1593 447 1599 453
rect 1605 447 1608 453
rect -84 444 1608 447
rect -84 441 -72 444
rect -84 435 -81 441
rect -75 435 -72 441
rect -84 429 -72 435
rect 1596 441 1608 444
rect 1596 435 1599 441
rect 1605 435 1608 441
rect -84 423 -81 429
rect -75 423 -72 429
rect 1596 429 1608 435
rect -84 417 -72 423
rect -84 411 -81 417
rect -75 411 -72 417
rect -84 405 -72 411
rect -84 399 -81 405
rect -75 399 -72 405
rect -84 393 -72 399
rect 1596 423 1599 429
rect 1605 423 1608 429
rect 1596 417 1608 423
rect 1596 411 1599 417
rect 1605 411 1608 417
rect 1596 405 1608 411
rect 1596 399 1599 405
rect 1605 399 1608 405
rect -84 387 -81 393
rect -75 387 -72 393
rect -84 381 -72 387
rect -84 375 -81 381
rect -75 375 -72 381
rect -84 369 -72 375
rect 1596 393 1608 399
rect 1596 387 1599 393
rect 1605 387 1608 393
rect 1596 381 1608 387
rect 1596 375 1599 381
rect 1605 375 1608 381
rect -84 363 -81 369
rect -75 363 -72 369
rect -84 360 -72 363
rect 1596 369 1608 375
rect 1596 363 1599 369
rect 1605 363 1608 369
rect 1596 360 1608 363
rect -84 357 1608 360
rect -84 351 -81 357
rect -75 351 -69 357
rect -63 351 -57 357
rect -51 351 -45 357
rect -39 351 -33 357
rect -27 351 -21 357
rect -15 351 -9 357
rect -3 351 3 357
rect 9 351 15 357
rect 21 351 27 357
rect 33 351 39 357
rect 45 351 51 357
rect 57 351 63 357
rect 69 351 75 357
rect 81 351 87 357
rect 93 351 99 357
rect 105 351 111 357
rect 117 351 123 357
rect 129 351 135 357
rect 141 351 147 357
rect 153 351 159 357
rect 165 351 171 357
rect 177 351 183 357
rect 189 351 195 357
rect 201 351 207 357
rect 213 351 219 357
rect 225 351 231 357
rect 237 351 243 357
rect 249 351 255 357
rect 261 351 267 357
rect 273 351 279 357
rect 285 351 291 357
rect 297 351 303 357
rect 309 351 315 357
rect 321 351 327 357
rect 333 351 339 357
rect 345 351 351 357
rect 357 351 363 357
rect 369 351 375 357
rect 381 351 387 357
rect 393 351 399 357
rect 405 351 411 357
rect 417 351 423 357
rect 429 351 435 357
rect 441 351 447 357
rect 453 351 459 357
rect 465 351 471 357
rect 477 351 483 357
rect 489 351 495 357
rect 501 351 507 357
rect 513 351 519 357
rect 525 351 531 357
rect 537 351 543 357
rect 549 351 555 357
rect 561 351 567 357
rect 573 351 579 357
rect 585 351 591 357
rect 597 351 603 357
rect 609 351 615 357
rect 621 351 627 357
rect 633 351 639 357
rect 645 351 651 357
rect 657 351 663 357
rect 669 351 675 357
rect 681 351 687 357
rect 693 351 699 357
rect 705 351 711 357
rect 717 351 723 357
rect 729 351 735 357
rect 741 351 747 357
rect 753 351 759 357
rect 765 351 771 357
rect 777 351 783 357
rect 789 351 795 357
rect 801 351 807 357
rect 813 351 819 357
rect 825 351 831 357
rect 837 351 843 357
rect 849 351 855 357
rect 861 351 867 357
rect 873 351 879 357
rect 885 351 891 357
rect 897 351 903 357
rect 909 351 915 357
rect 921 351 927 357
rect 933 351 939 357
rect 945 351 951 357
rect 957 351 963 357
rect 969 351 975 357
rect 981 351 987 357
rect 993 351 999 357
rect 1005 351 1011 357
rect 1017 351 1023 357
rect 1029 351 1035 357
rect 1041 351 1047 357
rect 1053 351 1059 357
rect 1065 351 1071 357
rect 1077 351 1083 357
rect 1089 351 1095 357
rect 1101 351 1107 357
rect 1113 351 1119 357
rect 1125 351 1131 357
rect 1137 351 1143 357
rect 1149 351 1155 357
rect 1161 351 1167 357
rect 1173 351 1179 357
rect 1185 351 1191 357
rect 1197 351 1203 357
rect 1209 351 1215 357
rect 1221 351 1227 357
rect 1233 351 1239 357
rect 1245 351 1251 357
rect 1257 351 1263 357
rect 1269 351 1275 357
rect 1281 351 1287 357
rect 1293 351 1299 357
rect 1305 351 1311 357
rect 1317 351 1323 357
rect 1329 351 1335 357
rect 1341 351 1347 357
rect 1353 351 1359 357
rect 1365 351 1371 357
rect 1377 351 1383 357
rect 1389 351 1395 357
rect 1401 351 1407 357
rect 1413 351 1419 357
rect 1425 351 1431 357
rect 1437 351 1443 357
rect 1449 351 1455 357
rect 1461 351 1467 357
rect 1473 351 1479 357
rect 1485 351 1491 357
rect 1497 351 1503 357
rect 1509 351 1515 357
rect 1521 351 1527 357
rect 1533 351 1539 357
rect 1545 351 1551 357
rect 1557 351 1563 357
rect 1569 351 1575 357
rect 1581 351 1587 357
rect 1593 351 1599 357
rect 1605 351 1608 357
rect -84 348 1608 351
<< mvnsubdiff >>
rect -60 501 1584 504
rect -60 495 -57 501
rect -51 495 -45 501
rect -39 495 -33 501
rect -27 495 -21 501
rect -15 495 -9 501
rect -3 495 3 501
rect 9 495 15 501
rect 21 495 27 501
rect 33 495 39 501
rect 45 495 51 501
rect 57 495 63 501
rect 69 495 75 501
rect 81 495 87 501
rect 93 495 99 501
rect 105 495 111 501
rect 117 495 123 501
rect 129 495 135 501
rect 141 495 147 501
rect 153 495 159 501
rect 165 495 171 501
rect 177 495 183 501
rect 189 495 195 501
rect 201 495 207 501
rect 213 495 219 501
rect 225 495 231 501
rect 237 495 243 501
rect 249 495 255 501
rect 261 495 267 501
rect 273 495 279 501
rect 285 495 291 501
rect 297 495 303 501
rect 309 495 315 501
rect 321 495 327 501
rect 333 495 339 501
rect 345 495 351 501
rect 357 495 363 501
rect 369 495 375 501
rect 381 495 387 501
rect 393 495 399 501
rect 405 495 411 501
rect 417 495 423 501
rect 429 495 435 501
rect 441 495 447 501
rect 453 495 459 501
rect 465 495 471 501
rect 477 495 483 501
rect 489 495 495 501
rect 501 495 507 501
rect 513 495 519 501
rect 525 495 531 501
rect 537 495 543 501
rect 549 495 555 501
rect 561 495 567 501
rect 573 495 579 501
rect 585 495 591 501
rect 597 495 603 501
rect 609 495 615 501
rect 621 495 627 501
rect 633 495 639 501
rect 645 495 651 501
rect 657 495 663 501
rect 669 495 675 501
rect 681 495 687 501
rect 693 495 699 501
rect 705 495 711 501
rect 717 495 723 501
rect 729 495 735 501
rect 741 495 747 501
rect 753 495 759 501
rect 765 495 771 501
rect 777 495 783 501
rect 789 495 795 501
rect 801 495 807 501
rect 813 495 819 501
rect 825 495 831 501
rect 837 495 843 501
rect 849 495 855 501
rect 861 495 867 501
rect 873 495 879 501
rect 885 495 891 501
rect 897 495 903 501
rect 909 495 915 501
rect 921 495 927 501
rect 933 495 939 501
rect 945 495 951 501
rect 957 495 963 501
rect 969 495 975 501
rect 981 495 987 501
rect 993 495 999 501
rect 1005 495 1011 501
rect 1017 495 1023 501
rect 1029 495 1035 501
rect 1041 495 1047 501
rect 1053 495 1059 501
rect 1065 495 1071 501
rect 1077 495 1083 501
rect 1089 495 1095 501
rect 1101 495 1107 501
rect 1113 495 1119 501
rect 1125 495 1131 501
rect 1137 495 1143 501
rect 1149 495 1155 501
rect 1161 495 1167 501
rect 1173 495 1179 501
rect 1185 495 1191 501
rect 1197 495 1203 501
rect 1209 495 1215 501
rect 1221 495 1227 501
rect 1233 495 1239 501
rect 1245 495 1251 501
rect 1257 495 1263 501
rect 1269 495 1275 501
rect 1281 495 1287 501
rect 1293 495 1299 501
rect 1305 495 1311 501
rect 1317 495 1323 501
rect 1329 495 1335 501
rect 1341 495 1347 501
rect 1353 495 1359 501
rect 1365 495 1371 501
rect 1377 495 1383 501
rect 1389 495 1395 501
rect 1401 495 1407 501
rect 1413 495 1419 501
rect 1425 495 1431 501
rect 1437 495 1443 501
rect 1449 495 1455 501
rect 1461 495 1467 501
rect 1473 495 1479 501
rect 1485 495 1491 501
rect 1497 495 1503 501
rect 1509 495 1515 501
rect 1521 495 1527 501
rect 1533 495 1539 501
rect 1545 495 1551 501
rect 1557 495 1563 501
rect 1569 495 1575 501
rect 1581 495 1584 501
rect -60 492 1584 495
<< psubdiffcont >>
rect -105 615 -99 621
rect -93 615 -87 621
rect -81 615 -75 621
rect -69 615 -63 621
rect -57 615 -51 621
rect -45 615 -39 621
rect -33 615 -27 621
rect -21 615 -15 621
rect -9 615 -3 621
rect 3 615 9 621
rect 15 615 21 621
rect 27 615 33 621
rect 39 615 45 621
rect 51 615 57 621
rect 63 615 69 621
rect 75 615 81 621
rect 87 615 93 621
rect 99 615 105 621
rect 111 615 117 621
rect 123 615 129 621
rect 135 615 141 621
rect 147 615 153 621
rect 159 615 165 621
rect 171 615 177 621
rect 183 615 189 621
rect 195 615 201 621
rect 207 615 213 621
rect 219 615 225 621
rect 231 615 237 621
rect 243 615 249 621
rect 255 615 261 621
rect 267 615 273 621
rect 279 615 285 621
rect 291 615 297 621
rect 303 615 309 621
rect 315 615 321 621
rect 327 615 333 621
rect 339 615 345 621
rect 351 615 357 621
rect 363 615 369 621
rect 375 615 381 621
rect 387 615 393 621
rect 399 615 405 621
rect 411 615 417 621
rect 423 615 429 621
rect 435 615 441 621
rect 447 615 453 621
rect 459 615 465 621
rect 471 615 477 621
rect 483 615 489 621
rect 495 615 501 621
rect 507 615 513 621
rect 519 615 525 621
rect 531 615 537 621
rect 543 615 549 621
rect 555 615 561 621
rect 567 615 573 621
rect 579 615 585 621
rect 591 615 597 621
rect 603 615 609 621
rect 615 615 621 621
rect 627 615 633 621
rect 639 615 645 621
rect 651 615 657 621
rect 663 615 669 621
rect 675 615 681 621
rect 687 615 693 621
rect 699 615 705 621
rect 711 615 717 621
rect 723 615 729 621
rect 735 615 741 621
rect 747 615 753 621
rect 759 615 765 621
rect 771 615 777 621
rect 783 615 789 621
rect 795 615 801 621
rect 807 615 813 621
rect 819 615 825 621
rect 831 615 837 621
rect 843 615 849 621
rect 855 615 861 621
rect 867 615 873 621
rect 879 615 885 621
rect 891 615 897 621
rect 903 615 909 621
rect 915 615 921 621
rect 927 615 933 621
rect 939 615 945 621
rect 951 615 957 621
rect 963 615 969 621
rect 975 615 981 621
rect 987 615 993 621
rect 999 615 1005 621
rect 1011 615 1017 621
rect 1023 615 1029 621
rect 1035 615 1041 621
rect 1047 615 1053 621
rect 1059 615 1065 621
rect 1071 615 1077 621
rect 1083 615 1089 621
rect 1095 615 1101 621
rect 1107 615 1113 621
rect 1119 615 1125 621
rect 1131 615 1137 621
rect 1143 615 1149 621
rect 1155 615 1161 621
rect 1167 615 1173 621
rect 1179 615 1185 621
rect 1191 615 1197 621
rect 1203 615 1209 621
rect 1215 615 1221 621
rect 1227 615 1233 621
rect 1239 615 1245 621
rect 1251 615 1257 621
rect 1263 615 1269 621
rect 1275 615 1281 621
rect 1287 615 1293 621
rect 1299 615 1305 621
rect 1311 615 1317 621
rect 1323 615 1329 621
rect 1335 615 1341 621
rect 1347 615 1353 621
rect 1359 615 1365 621
rect 1371 615 1377 621
rect 1383 615 1389 621
rect 1395 615 1401 621
rect 1407 615 1413 621
rect 1419 615 1425 621
rect 1431 615 1437 621
rect 1443 615 1449 621
rect 1455 615 1461 621
rect 1467 615 1473 621
rect 1479 615 1485 621
rect 1491 615 1497 621
rect 1503 615 1509 621
rect 1515 615 1521 621
rect 1527 615 1533 621
rect 1539 615 1545 621
rect 1551 615 1557 621
rect 1563 615 1569 621
rect 1575 615 1581 621
rect 1587 615 1593 621
rect 1599 615 1605 621
rect 1611 615 1617 621
rect 1623 615 1629 621
rect -105 603 -99 609
rect 1623 603 1629 609
rect -105 591 -99 597
rect -105 579 -99 585
rect -105 567 -99 573
rect -105 555 -99 561
rect -105 543 -99 549
rect -105 531 -99 537
rect -105 519 -99 525
rect -105 507 -99 513
rect -105 495 -99 501
rect 1623 591 1629 597
rect 1623 579 1629 585
rect 1623 567 1629 573
rect 1623 555 1629 561
rect 1623 543 1629 549
rect 1623 531 1629 537
rect 1623 519 1629 525
rect 1623 507 1629 513
rect 1623 495 1629 501
rect -105 483 -99 489
rect 1623 483 1629 489
rect -105 471 -99 477
rect -93 471 -87 477
rect -81 471 -75 477
rect -69 471 -63 477
rect -57 471 -51 477
rect -45 471 -39 477
rect -33 471 -27 477
rect -21 471 -15 477
rect -9 471 -3 477
rect 3 471 9 477
rect 15 471 21 477
rect 27 471 33 477
rect 39 471 45 477
rect 51 471 57 477
rect 63 471 69 477
rect 75 471 81 477
rect 87 471 93 477
rect 99 471 105 477
rect 111 471 117 477
rect 123 471 129 477
rect 135 471 141 477
rect 147 471 153 477
rect 159 471 165 477
rect 171 471 177 477
rect 183 471 189 477
rect 195 471 201 477
rect 207 471 213 477
rect 219 471 225 477
rect 231 471 237 477
rect 243 471 249 477
rect 255 471 261 477
rect 267 471 273 477
rect 279 471 285 477
rect 291 471 297 477
rect 303 471 309 477
rect 315 471 321 477
rect 327 471 333 477
rect 339 471 345 477
rect 351 471 357 477
rect 363 471 369 477
rect 375 471 381 477
rect 387 471 393 477
rect 399 471 405 477
rect 411 471 417 477
rect 423 471 429 477
rect 435 471 441 477
rect 447 471 453 477
rect 459 471 465 477
rect 471 471 477 477
rect 483 471 489 477
rect 495 471 501 477
rect 507 471 513 477
rect 519 471 525 477
rect 531 471 537 477
rect 543 471 549 477
rect 555 471 561 477
rect 567 471 573 477
rect 579 471 585 477
rect 591 471 597 477
rect 603 471 609 477
rect 615 471 621 477
rect 627 471 633 477
rect 639 471 645 477
rect 651 471 657 477
rect 663 471 669 477
rect 675 471 681 477
rect 687 471 693 477
rect 699 471 705 477
rect 711 471 717 477
rect 723 471 729 477
rect 735 471 741 477
rect 747 471 753 477
rect 759 471 765 477
rect 771 471 777 477
rect 783 471 789 477
rect 795 471 801 477
rect 807 471 813 477
rect 819 471 825 477
rect 831 471 837 477
rect 843 471 849 477
rect 855 471 861 477
rect 867 471 873 477
rect 879 471 885 477
rect 891 471 897 477
rect 903 471 909 477
rect 915 471 921 477
rect 927 471 933 477
rect 939 471 945 477
rect 951 471 957 477
rect 963 471 969 477
rect 975 471 981 477
rect 987 471 993 477
rect 999 471 1005 477
rect 1011 471 1017 477
rect 1023 471 1029 477
rect 1035 471 1041 477
rect 1047 471 1053 477
rect 1059 471 1065 477
rect 1071 471 1077 477
rect 1083 471 1089 477
rect 1095 471 1101 477
rect 1107 471 1113 477
rect 1119 471 1125 477
rect 1131 471 1137 477
rect 1143 471 1149 477
rect 1155 471 1161 477
rect 1167 471 1173 477
rect 1179 471 1185 477
rect 1191 471 1197 477
rect 1203 471 1209 477
rect 1215 471 1221 477
rect 1227 471 1233 477
rect 1239 471 1245 477
rect 1251 471 1257 477
rect 1263 471 1269 477
rect 1275 471 1281 477
rect 1287 471 1293 477
rect 1299 471 1305 477
rect 1311 471 1317 477
rect 1323 471 1329 477
rect 1335 471 1341 477
rect 1347 471 1353 477
rect 1359 471 1365 477
rect 1371 471 1377 477
rect 1383 471 1389 477
rect 1395 471 1401 477
rect 1407 471 1413 477
rect 1419 471 1425 477
rect 1431 471 1437 477
rect 1443 471 1449 477
rect 1455 471 1461 477
rect 1467 471 1473 477
rect 1479 471 1485 477
rect 1491 471 1497 477
rect 1503 471 1509 477
rect 1515 471 1521 477
rect 1527 471 1533 477
rect 1539 471 1545 477
rect 1551 471 1557 477
rect 1563 471 1569 477
rect 1575 471 1581 477
rect 1587 471 1593 477
rect 1599 471 1605 477
rect 1611 471 1617 477
rect 1623 471 1629 477
rect -105 459 -99 465
rect 1623 459 1629 465
rect -105 447 -99 453
rect -105 435 -99 441
rect -105 423 -99 429
rect -105 411 -99 417
rect -105 399 -99 405
rect -105 387 -99 393
rect -105 375 -99 381
rect -105 363 -99 369
rect -105 351 -99 357
rect 1623 447 1629 453
rect 1623 435 1629 441
rect 1623 423 1629 429
rect 1623 411 1629 417
rect 1623 399 1629 405
rect 1623 387 1629 393
rect 1623 375 1629 381
rect 1623 363 1629 369
rect 1623 351 1629 357
rect -105 339 -99 345
rect 1623 339 1629 345
rect -105 327 -99 333
rect -93 327 -87 333
rect -81 327 -75 333
rect -69 327 -63 333
rect -57 327 -51 333
rect -45 327 -39 333
rect -33 327 -27 333
rect -21 327 -15 333
rect -9 327 -3 333
rect 3 327 9 333
rect 15 327 21 333
rect 27 327 33 333
rect 39 327 45 333
rect 51 327 57 333
rect 63 327 69 333
rect 75 327 81 333
rect 87 327 93 333
rect 99 327 105 333
rect 111 327 117 333
rect 123 327 129 333
rect 135 327 141 333
rect 147 327 153 333
rect 159 327 165 333
rect 171 327 177 333
rect 183 327 189 333
rect 195 327 201 333
rect 207 327 213 333
rect 219 327 225 333
rect 231 327 237 333
rect 243 327 249 333
rect 255 327 261 333
rect 267 327 273 333
rect 279 327 285 333
rect 291 327 297 333
rect 303 327 309 333
rect 315 327 321 333
rect 327 327 333 333
rect 339 327 345 333
rect 351 327 357 333
rect 363 327 369 333
rect 375 327 381 333
rect 387 327 393 333
rect 399 327 405 333
rect 411 327 417 333
rect 423 327 429 333
rect 435 327 441 333
rect 447 327 453 333
rect 459 327 465 333
rect 471 327 477 333
rect 483 327 489 333
rect 495 327 501 333
rect 507 327 513 333
rect 519 327 525 333
rect 531 327 537 333
rect 543 327 549 333
rect 555 327 561 333
rect 567 327 573 333
rect 579 327 585 333
rect 591 327 597 333
rect 603 327 609 333
rect 615 327 621 333
rect 627 327 633 333
rect 639 327 645 333
rect 651 327 657 333
rect 663 327 669 333
rect 675 327 681 333
rect 687 327 693 333
rect 699 327 705 333
rect 711 327 717 333
rect 723 327 729 333
rect 735 327 741 333
rect 747 327 753 333
rect 759 327 765 333
rect 771 327 777 333
rect 783 327 789 333
rect 795 327 801 333
rect 807 327 813 333
rect 819 327 825 333
rect 831 327 837 333
rect 843 327 849 333
rect 855 327 861 333
rect 867 327 873 333
rect 879 327 885 333
rect 891 327 897 333
rect 903 327 909 333
rect 915 327 921 333
rect 927 327 933 333
rect 939 327 945 333
rect 951 327 957 333
rect 963 327 969 333
rect 975 327 981 333
rect 987 327 993 333
rect 999 327 1005 333
rect 1011 327 1017 333
rect 1023 327 1029 333
rect 1035 327 1041 333
rect 1047 327 1053 333
rect 1059 327 1065 333
rect 1071 327 1077 333
rect 1083 327 1089 333
rect 1095 327 1101 333
rect 1107 327 1113 333
rect 1119 327 1125 333
rect 1131 327 1137 333
rect 1143 327 1149 333
rect 1155 327 1161 333
rect 1167 327 1173 333
rect 1179 327 1185 333
rect 1191 327 1197 333
rect 1203 327 1209 333
rect 1215 327 1221 333
rect 1227 327 1233 333
rect 1239 327 1245 333
rect 1251 327 1257 333
rect 1263 327 1269 333
rect 1275 327 1281 333
rect 1287 327 1293 333
rect 1299 327 1305 333
rect 1311 327 1317 333
rect 1323 327 1329 333
rect 1335 327 1341 333
rect 1347 327 1353 333
rect 1359 327 1365 333
rect 1371 327 1377 333
rect 1383 327 1389 333
rect 1395 327 1401 333
rect 1407 327 1413 333
rect 1419 327 1425 333
rect 1431 327 1437 333
rect 1443 327 1449 333
rect 1455 327 1461 333
rect 1467 327 1473 333
rect 1479 327 1485 333
rect 1491 327 1497 333
rect 1503 327 1509 333
rect 1515 327 1521 333
rect 1527 327 1533 333
rect 1539 327 1545 333
rect 1551 327 1557 333
rect 1563 327 1569 333
rect 1575 327 1581 333
rect 1587 327 1593 333
rect 1599 327 1605 333
rect 1611 327 1617 333
rect 1623 327 1629 333
rect -105 315 -99 321
rect -105 303 -99 309
rect -105 291 -99 297
rect -105 279 -99 285
rect -105 267 -99 273
rect -105 255 -99 261
rect -105 243 -99 249
rect -105 231 -99 237
rect -105 219 -99 225
rect -105 207 -99 213
rect -105 195 -99 201
rect -105 183 -99 189
rect -105 171 -99 177
rect -105 159 -99 165
rect -105 147 -99 153
rect -105 135 -99 141
rect -105 123 -99 129
rect -105 111 -99 117
rect -105 99 -99 105
rect 1623 315 1629 321
rect 1623 303 1629 309
rect 1623 291 1629 297
rect 1623 279 1629 285
rect 1623 267 1629 273
rect 1623 255 1629 261
rect 1623 243 1629 249
rect 1623 231 1629 237
rect 1623 219 1629 225
rect 1623 207 1629 213
rect 1623 195 1629 201
rect 1623 183 1629 189
rect 1623 171 1629 177
rect 1623 159 1629 165
rect 1623 147 1629 153
rect 1623 135 1629 141
rect 1623 123 1629 129
rect 1623 111 1629 117
rect 1623 99 1629 105
rect -105 87 -99 93
rect -93 87 -87 93
rect -81 87 -75 93
rect -69 87 -63 93
rect -57 87 -51 93
rect -45 87 -39 93
rect -33 87 -27 93
rect -21 87 -15 93
rect -9 87 -3 93
rect 3 87 9 93
rect 15 87 21 93
rect 27 87 33 93
rect 39 87 45 93
rect 51 87 57 93
rect 63 87 69 93
rect 75 87 81 93
rect 87 87 93 93
rect 99 87 105 93
rect 111 87 117 93
rect 123 87 129 93
rect 135 87 141 93
rect 147 87 153 93
rect 159 87 165 93
rect 171 87 177 93
rect 183 87 189 93
rect 195 87 201 93
rect 207 87 213 93
rect 219 87 225 93
rect 231 87 237 93
rect 243 87 249 93
rect 255 87 261 93
rect 267 87 273 93
rect 279 87 285 93
rect 291 87 297 93
rect 303 87 309 93
rect 315 87 321 93
rect 327 87 333 93
rect 339 87 345 93
rect 351 87 357 93
rect 363 87 369 93
rect 375 87 381 93
rect 387 87 393 93
rect 399 87 405 93
rect 411 87 417 93
rect 423 87 429 93
rect 435 87 441 93
rect 447 87 453 93
rect 459 87 465 93
rect 471 87 477 93
rect 483 87 489 93
rect 495 87 501 93
rect 507 87 513 93
rect 519 87 525 93
rect 531 87 537 93
rect 543 87 549 93
rect 555 87 561 93
rect 567 87 573 93
rect 579 87 585 93
rect 591 87 597 93
rect 603 87 609 93
rect 615 87 621 93
rect 627 87 633 93
rect 639 87 645 93
rect 651 87 657 93
rect 663 87 669 93
rect 675 87 681 93
rect 687 87 693 93
rect 699 87 705 93
rect 711 87 717 93
rect 723 87 729 93
rect 735 87 741 93
rect 747 87 753 93
rect 759 87 765 93
rect 771 87 777 93
rect 783 87 789 93
rect 795 87 801 93
rect 807 87 813 93
rect 819 87 825 93
rect 831 87 837 93
rect 843 87 849 93
rect 855 87 861 93
rect 867 87 873 93
rect 879 87 885 93
rect 891 87 897 93
rect 903 87 909 93
rect 915 87 921 93
rect 927 87 933 93
rect 939 87 945 93
rect 951 87 957 93
rect 963 87 969 93
rect 975 87 981 93
rect 987 87 993 93
rect 999 87 1005 93
rect 1011 87 1017 93
rect 1023 87 1029 93
rect 1035 87 1041 93
rect 1047 87 1053 93
rect 1059 87 1065 93
rect 1071 87 1077 93
rect 1083 87 1089 93
rect 1095 87 1101 93
rect 1107 87 1113 93
rect 1119 87 1125 93
rect 1131 87 1137 93
rect 1143 87 1149 93
rect 1155 87 1161 93
rect 1167 87 1173 93
rect 1179 87 1185 93
rect 1191 87 1197 93
rect 1203 87 1209 93
rect 1215 87 1221 93
rect 1227 87 1233 93
rect 1239 87 1245 93
rect 1251 87 1257 93
rect 1263 87 1269 93
rect 1275 87 1281 93
rect 1287 87 1293 93
rect 1299 87 1305 93
rect 1311 87 1317 93
rect 1323 87 1329 93
rect 1335 87 1341 93
rect 1347 87 1353 93
rect 1359 87 1365 93
rect 1371 87 1377 93
rect 1383 87 1389 93
rect 1395 87 1401 93
rect 1407 87 1413 93
rect 1419 87 1425 93
rect 1431 87 1437 93
rect 1443 87 1449 93
rect 1455 87 1461 93
rect 1467 87 1473 93
rect 1479 87 1485 93
rect 1491 87 1497 93
rect 1503 87 1509 93
rect 1515 87 1521 93
rect 1527 87 1533 93
rect 1539 87 1545 93
rect 1551 87 1557 93
rect 1563 87 1569 93
rect 1575 87 1581 93
rect 1587 87 1593 93
rect 1599 87 1605 93
rect 1611 87 1617 93
rect 1623 87 1629 93
rect -105 75 -99 81
rect 1623 75 1629 81
rect -105 63 -99 69
rect -105 51 -99 57
rect 1623 63 1629 69
rect 1623 51 1629 57
rect -105 39 -99 45
rect -105 27 -99 33
rect -105 15 -99 21
rect 1623 39 1629 45
rect 1623 27 1629 33
rect 1623 15 1629 21
rect -105 3 -99 9
rect 1623 3 1629 9
rect -105 -9 -99 -3
rect -93 -9 -87 -3
rect -81 -9 -75 -3
rect -69 -9 -63 -3
rect -57 -9 -51 -3
rect -45 -9 -39 -3
rect -33 -9 -27 -3
rect -21 -9 -15 -3
rect -9 -9 -3 -3
rect 3 -9 9 -3
rect 15 -9 21 -3
rect 27 -9 33 -3
rect 39 -9 45 -3
rect 51 -9 57 -3
rect 63 -9 69 -3
rect 75 -9 81 -3
rect 87 -9 93 -3
rect 99 -9 105 -3
rect 111 -9 117 -3
rect 123 -9 129 -3
rect 135 -9 141 -3
rect 147 -9 153 -3
rect 159 -9 165 -3
rect 171 -9 177 -3
rect 183 -9 189 -3
rect 195 -9 201 -3
rect 207 -9 213 -3
rect 219 -9 225 -3
rect 231 -9 237 -3
rect 243 -9 249 -3
rect 255 -9 261 -3
rect 267 -9 273 -3
rect 279 -9 285 -3
rect 291 -9 297 -3
rect 303 -9 309 -3
rect 315 -9 321 -3
rect 327 -9 333 -3
rect 339 -9 345 -3
rect 351 -9 357 -3
rect 363 -9 369 -3
rect 375 -9 381 -3
rect 387 -9 393 -3
rect 399 -9 405 -3
rect 411 -9 417 -3
rect 423 -9 429 -3
rect 435 -9 441 -3
rect 447 -9 453 -3
rect 459 -9 465 -3
rect 471 -9 477 -3
rect 483 -9 489 -3
rect 495 -9 501 -3
rect 507 -9 513 -3
rect 519 -9 525 -3
rect 531 -9 537 -3
rect 543 -9 549 -3
rect 555 -9 561 -3
rect 567 -9 573 -3
rect 579 -9 585 -3
rect 591 -9 597 -3
rect 603 -9 609 -3
rect 615 -9 621 -3
rect 627 -9 633 -3
rect 639 -9 645 -3
rect 651 -9 657 -3
rect 663 -9 669 -3
rect 675 -9 681 -3
rect 687 -9 693 -3
rect 699 -9 705 -3
rect 711 -9 717 -3
rect 723 -9 729 -3
rect 735 -9 741 -3
rect 747 -9 753 -3
rect 759 -9 765 -3
rect 771 -9 777 -3
rect 783 -9 789 -3
rect 795 -9 801 -3
rect 807 -9 813 -3
rect 819 -9 825 -3
rect 831 -9 837 -3
rect 843 -9 849 -3
rect 855 -9 861 -3
rect 867 -9 873 -3
rect 879 -9 885 -3
rect 891 -9 897 -3
rect 903 -9 909 -3
rect 915 -9 921 -3
rect 927 -9 933 -3
rect 939 -9 945 -3
rect 951 -9 957 -3
rect 963 -9 969 -3
rect 975 -9 981 -3
rect 987 -9 993 -3
rect 999 -9 1005 -3
rect 1011 -9 1017 -3
rect 1023 -9 1029 -3
rect 1035 -9 1041 -3
rect 1047 -9 1053 -3
rect 1059 -9 1065 -3
rect 1071 -9 1077 -3
rect 1083 -9 1089 -3
rect 1095 -9 1101 -3
rect 1107 -9 1113 -3
rect 1119 -9 1125 -3
rect 1131 -9 1137 -3
rect 1143 -9 1149 -3
rect 1155 -9 1161 -3
rect 1167 -9 1173 -3
rect 1179 -9 1185 -3
rect 1191 -9 1197 -3
rect 1203 -9 1209 -3
rect 1215 -9 1221 -3
rect 1227 -9 1233 -3
rect 1239 -9 1245 -3
rect 1251 -9 1257 -3
rect 1263 -9 1269 -3
rect 1275 -9 1281 -3
rect 1287 -9 1293 -3
rect 1299 -9 1305 -3
rect 1311 -9 1317 -3
rect 1323 -9 1329 -3
rect 1335 -9 1341 -3
rect 1347 -9 1353 -3
rect 1359 -9 1365 -3
rect 1371 -9 1377 -3
rect 1383 -9 1389 -3
rect 1395 -9 1401 -3
rect 1407 -9 1413 -3
rect 1419 -9 1425 -3
rect 1431 -9 1437 -3
rect 1443 -9 1449 -3
rect 1455 -9 1461 -3
rect 1467 -9 1473 -3
rect 1479 -9 1485 -3
rect 1491 -9 1497 -3
rect 1503 -9 1509 -3
rect 1515 -9 1521 -3
rect 1527 -9 1533 -3
rect 1539 -9 1545 -3
rect 1551 -9 1557 -3
rect 1563 -9 1569 -3
rect 1575 -9 1581 -3
rect 1587 -9 1593 -3
rect 1599 -9 1605 -3
rect 1611 -9 1617 -3
rect 1623 -9 1629 -3
rect -105 -21 -99 -15
rect -105 -33 -99 -27
rect -105 -45 -99 -39
rect -105 -57 -99 -51
rect -105 -69 -99 -63
rect -105 -81 -99 -75
rect -105 -93 -99 -87
rect -105 -105 -99 -99
rect -105 -117 -99 -111
rect -105 -129 -99 -123
rect -105 -141 -99 -135
rect -105 -153 -99 -147
rect -105 -165 -99 -159
rect -105 -177 -99 -171
rect -105 -189 -99 -183
rect 1623 -21 1629 -15
rect 1623 -33 1629 -27
rect 1623 -45 1629 -39
rect 1623 -57 1629 -51
rect 1623 -69 1629 -63
rect 1623 -81 1629 -75
rect 1623 -93 1629 -87
rect 1623 -105 1629 -99
rect 1623 -117 1629 -111
rect 1623 -129 1629 -123
rect 1623 -141 1629 -135
rect 1623 -153 1629 -147
rect 1623 -165 1629 -159
rect 1623 -177 1629 -171
rect 1623 -189 1629 -183
rect -105 -201 -99 -195
rect -93 -201 -87 -195
rect -81 -201 -75 -195
rect -69 -201 -63 -195
rect -57 -201 -51 -195
rect -45 -201 -39 -195
rect -33 -201 -27 -195
rect -21 -201 -15 -195
rect -9 -201 -3 -195
rect 3 -201 9 -195
rect 15 -201 21 -195
rect 27 -201 33 -195
rect 39 -201 45 -195
rect 51 -201 57 -195
rect 63 -201 69 -195
rect 75 -201 81 -195
rect 87 -201 93 -195
rect 99 -201 105 -195
rect 111 -201 117 -195
rect 123 -201 129 -195
rect 135 -201 141 -195
rect 147 -201 153 -195
rect 159 -201 165 -195
rect 171 -201 177 -195
rect 183 -201 189 -195
rect 195 -201 201 -195
rect 207 -201 213 -195
rect 219 -201 225 -195
rect 231 -201 237 -195
rect 243 -201 249 -195
rect 255 -201 261 -195
rect 267 -201 273 -195
rect 279 -201 285 -195
rect 291 -201 297 -195
rect 303 -201 309 -195
rect 315 -201 321 -195
rect 327 -201 333 -195
rect 339 -201 345 -195
rect 351 -201 357 -195
rect 363 -201 369 -195
rect 375 -201 381 -195
rect 387 -201 393 -195
rect 399 -201 405 -195
rect 411 -201 417 -195
rect 423 -201 429 -195
rect 435 -201 441 -195
rect 447 -201 453 -195
rect 459 -201 465 -195
rect 471 -201 477 -195
rect 483 -201 489 -195
rect 495 -201 501 -195
rect 507 -201 513 -195
rect 519 -201 525 -195
rect 531 -201 537 -195
rect 543 -201 549 -195
rect 555 -201 561 -195
rect 567 -201 573 -195
rect 579 -201 585 -195
rect 591 -201 597 -195
rect 603 -201 609 -195
rect 615 -201 621 -195
rect 627 -201 633 -195
rect 639 -201 645 -195
rect 651 -201 657 -195
rect 663 -201 669 -195
rect 675 -201 681 -195
rect 687 -201 693 -195
rect 699 -201 705 -195
rect 711 -201 717 -195
rect 723 -201 729 -195
rect 735 -201 741 -195
rect 747 -201 753 -195
rect 759 -201 765 -195
rect 771 -201 777 -195
rect 783 -201 789 -195
rect 795 -201 801 -195
rect 807 -201 813 -195
rect 819 -201 825 -195
rect 831 -201 837 -195
rect 843 -201 849 -195
rect 855 -201 861 -195
rect 867 -201 873 -195
rect 879 -201 885 -195
rect 891 -201 897 -195
rect 903 -201 909 -195
rect 915 -201 921 -195
rect 927 -201 933 -195
rect 939 -201 945 -195
rect 951 -201 957 -195
rect 963 -201 969 -195
rect 975 -201 981 -195
rect 987 -201 993 -195
rect 999 -201 1005 -195
rect 1011 -201 1017 -195
rect 1023 -201 1029 -195
rect 1035 -201 1041 -195
rect 1047 -201 1053 -195
rect 1059 -201 1065 -195
rect 1071 -201 1077 -195
rect 1083 -201 1089 -195
rect 1095 -201 1101 -195
rect 1107 -201 1113 -195
rect 1119 -201 1125 -195
rect 1131 -201 1137 -195
rect 1143 -201 1149 -195
rect 1155 -201 1161 -195
rect 1167 -201 1173 -195
rect 1179 -201 1185 -195
rect 1191 -201 1197 -195
rect 1203 -201 1209 -195
rect 1215 -201 1221 -195
rect 1227 -201 1233 -195
rect 1239 -201 1245 -195
rect 1251 -201 1257 -195
rect 1263 -201 1269 -195
rect 1275 -201 1281 -195
rect 1287 -201 1293 -195
rect 1299 -201 1305 -195
rect 1311 -201 1317 -195
rect 1323 -201 1329 -195
rect 1335 -201 1341 -195
rect 1347 -201 1353 -195
rect 1359 -201 1365 -195
rect 1371 -201 1377 -195
rect 1383 -201 1389 -195
rect 1395 -201 1401 -195
rect 1407 -201 1413 -195
rect 1419 -201 1425 -195
rect 1431 -201 1437 -195
rect 1443 -201 1449 -195
rect 1455 -201 1461 -195
rect 1563 -201 1569 -195
rect 1575 -201 1581 -195
rect 1587 -201 1593 -195
rect 1599 -201 1605 -195
rect 1611 -201 1617 -195
rect 1623 -201 1629 -195
<< nsubdiffcont >>
rect -81 591 -75 597
rect -69 591 -63 597
rect -57 591 -51 597
rect -45 591 -39 597
rect -33 591 -27 597
rect -21 591 -15 597
rect -9 591 -3 597
rect 3 591 9 597
rect 15 591 21 597
rect 27 591 33 597
rect 39 591 45 597
rect 51 591 57 597
rect 63 591 69 597
rect 75 591 81 597
rect 87 591 93 597
rect 99 591 105 597
rect 111 591 117 597
rect 123 591 129 597
rect 135 591 141 597
rect 147 591 153 597
rect 159 591 165 597
rect 171 591 177 597
rect 183 591 189 597
rect 195 591 201 597
rect 207 591 213 597
rect 219 591 225 597
rect 231 591 237 597
rect 243 591 249 597
rect 255 591 261 597
rect 267 591 273 597
rect 279 591 285 597
rect 291 591 297 597
rect 303 591 309 597
rect 315 591 321 597
rect 327 591 333 597
rect 339 591 345 597
rect 351 591 357 597
rect 363 591 369 597
rect 375 591 381 597
rect 387 591 393 597
rect 399 591 405 597
rect 411 591 417 597
rect 423 591 429 597
rect 435 591 441 597
rect 447 591 453 597
rect 459 591 465 597
rect 471 591 477 597
rect 483 591 489 597
rect 495 591 501 597
rect 507 591 513 597
rect 519 591 525 597
rect 531 591 537 597
rect 543 591 549 597
rect 555 591 561 597
rect 567 591 573 597
rect 579 591 585 597
rect 591 591 597 597
rect 603 591 609 597
rect 615 591 621 597
rect 627 591 633 597
rect 639 591 645 597
rect 651 591 657 597
rect 663 591 669 597
rect 675 591 681 597
rect 687 591 693 597
rect 699 591 705 597
rect 711 591 717 597
rect 723 591 729 597
rect 735 591 741 597
rect 747 591 753 597
rect 759 591 765 597
rect 771 591 777 597
rect 783 591 789 597
rect 795 591 801 597
rect 807 591 813 597
rect 819 591 825 597
rect 831 591 837 597
rect 843 591 849 597
rect 855 591 861 597
rect 867 591 873 597
rect 879 591 885 597
rect 891 591 897 597
rect 903 591 909 597
rect 915 591 921 597
rect 927 591 933 597
rect 939 591 945 597
rect 951 591 957 597
rect 963 591 969 597
rect 975 591 981 597
rect 987 591 993 597
rect 999 591 1005 597
rect 1011 591 1017 597
rect 1023 591 1029 597
rect 1035 591 1041 597
rect 1047 591 1053 597
rect 1059 591 1065 597
rect 1071 591 1077 597
rect 1083 591 1089 597
rect 1095 591 1101 597
rect 1107 591 1113 597
rect 1119 591 1125 597
rect 1131 591 1137 597
rect 1143 591 1149 597
rect 1155 591 1161 597
rect 1167 591 1173 597
rect 1179 591 1185 597
rect 1191 591 1197 597
rect 1203 591 1209 597
rect 1215 591 1221 597
rect 1227 591 1233 597
rect 1239 591 1245 597
rect 1251 591 1257 597
rect 1263 591 1269 597
rect 1275 591 1281 597
rect 1287 591 1293 597
rect 1299 591 1305 597
rect 1311 591 1317 597
rect 1323 591 1329 597
rect 1335 591 1341 597
rect 1347 591 1353 597
rect 1359 591 1365 597
rect 1371 591 1377 597
rect 1383 591 1389 597
rect 1395 591 1401 597
rect 1407 591 1413 597
rect 1419 591 1425 597
rect 1431 591 1437 597
rect 1443 591 1449 597
rect 1455 591 1461 597
rect 1467 591 1473 597
rect 1479 591 1485 597
rect 1491 591 1497 597
rect 1503 591 1509 597
rect 1515 591 1521 597
rect 1527 591 1533 597
rect 1539 591 1545 597
rect 1551 591 1557 597
rect 1563 591 1569 597
rect 1575 591 1581 597
rect 1587 591 1593 597
rect 1599 591 1605 597
rect -81 579 -75 585
rect 1599 579 1605 585
rect -81 567 -75 573
rect -81 555 -75 561
rect 1599 567 1605 573
rect 1599 555 1605 561
rect -81 543 -75 549
rect -81 531 -75 537
rect -81 519 -75 525
rect 1599 543 1605 549
rect 1599 531 1605 537
rect 1599 519 1605 525
rect -81 507 -75 513
rect 1599 507 1605 513
rect -81 495 -75 501
rect -69 495 -63 501
rect 1587 495 1593 501
rect 1599 495 1605 501
rect -81 447 -75 453
rect -69 447 -63 453
rect -57 447 -51 453
rect -45 447 -39 453
rect -33 447 -27 453
rect -21 447 -15 453
rect -9 447 -3 453
rect 3 447 9 453
rect 15 447 21 453
rect 27 447 33 453
rect 39 447 45 453
rect 51 447 57 453
rect 63 447 69 453
rect 75 447 81 453
rect 87 447 93 453
rect 99 447 105 453
rect 111 447 117 453
rect 123 447 129 453
rect 135 447 141 453
rect 147 447 153 453
rect 159 447 165 453
rect 171 447 177 453
rect 183 447 189 453
rect 195 447 201 453
rect 207 447 213 453
rect 219 447 225 453
rect 231 447 237 453
rect 243 447 249 453
rect 255 447 261 453
rect 267 447 273 453
rect 279 447 285 453
rect 291 447 297 453
rect 303 447 309 453
rect 315 447 321 453
rect 327 447 333 453
rect 339 447 345 453
rect 351 447 357 453
rect 363 447 369 453
rect 375 447 381 453
rect 387 447 393 453
rect 399 447 405 453
rect 411 447 417 453
rect 423 447 429 453
rect 435 447 441 453
rect 447 447 453 453
rect 459 447 465 453
rect 471 447 477 453
rect 483 447 489 453
rect 495 447 501 453
rect 507 447 513 453
rect 519 447 525 453
rect 531 447 537 453
rect 543 447 549 453
rect 555 447 561 453
rect 567 447 573 453
rect 579 447 585 453
rect 591 447 597 453
rect 603 447 609 453
rect 615 447 621 453
rect 627 447 633 453
rect 639 447 645 453
rect 651 447 657 453
rect 663 447 669 453
rect 675 447 681 453
rect 687 447 693 453
rect 699 447 705 453
rect 711 447 717 453
rect 723 447 729 453
rect 735 447 741 453
rect 747 447 753 453
rect 759 447 765 453
rect 771 447 777 453
rect 783 447 789 453
rect 795 447 801 453
rect 807 447 813 453
rect 819 447 825 453
rect 831 447 837 453
rect 843 447 849 453
rect 855 447 861 453
rect 867 447 873 453
rect 879 447 885 453
rect 891 447 897 453
rect 903 447 909 453
rect 915 447 921 453
rect 927 447 933 453
rect 939 447 945 453
rect 951 447 957 453
rect 963 447 969 453
rect 975 447 981 453
rect 987 447 993 453
rect 999 447 1005 453
rect 1011 447 1017 453
rect 1023 447 1029 453
rect 1035 447 1041 453
rect 1047 447 1053 453
rect 1059 447 1065 453
rect 1071 447 1077 453
rect 1083 447 1089 453
rect 1095 447 1101 453
rect 1107 447 1113 453
rect 1119 447 1125 453
rect 1131 447 1137 453
rect 1143 447 1149 453
rect 1155 447 1161 453
rect 1167 447 1173 453
rect 1179 447 1185 453
rect 1191 447 1197 453
rect 1203 447 1209 453
rect 1215 447 1221 453
rect 1227 447 1233 453
rect 1239 447 1245 453
rect 1251 447 1257 453
rect 1263 447 1269 453
rect 1275 447 1281 453
rect 1287 447 1293 453
rect 1299 447 1305 453
rect 1311 447 1317 453
rect 1323 447 1329 453
rect 1335 447 1341 453
rect 1347 447 1353 453
rect 1359 447 1365 453
rect 1371 447 1377 453
rect 1383 447 1389 453
rect 1395 447 1401 453
rect 1407 447 1413 453
rect 1419 447 1425 453
rect 1431 447 1437 453
rect 1443 447 1449 453
rect 1455 447 1461 453
rect 1467 447 1473 453
rect 1479 447 1485 453
rect 1491 447 1497 453
rect 1503 447 1509 453
rect 1515 447 1521 453
rect 1527 447 1533 453
rect 1539 447 1545 453
rect 1551 447 1557 453
rect 1563 447 1569 453
rect 1575 447 1581 453
rect 1587 447 1593 453
rect 1599 447 1605 453
rect -81 435 -75 441
rect 1599 435 1605 441
rect -81 423 -75 429
rect -81 411 -75 417
rect -81 399 -75 405
rect 1599 423 1605 429
rect 1599 411 1605 417
rect 1599 399 1605 405
rect -81 387 -75 393
rect -81 375 -75 381
rect 1599 387 1605 393
rect 1599 375 1605 381
rect -81 363 -75 369
rect 1599 363 1605 369
rect -81 351 -75 357
rect -69 351 -63 357
rect -57 351 -51 357
rect -45 351 -39 357
rect -33 351 -27 357
rect -21 351 -15 357
rect -9 351 -3 357
rect 3 351 9 357
rect 15 351 21 357
rect 27 351 33 357
rect 39 351 45 357
rect 51 351 57 357
rect 63 351 69 357
rect 75 351 81 357
rect 87 351 93 357
rect 99 351 105 357
rect 111 351 117 357
rect 123 351 129 357
rect 135 351 141 357
rect 147 351 153 357
rect 159 351 165 357
rect 171 351 177 357
rect 183 351 189 357
rect 195 351 201 357
rect 207 351 213 357
rect 219 351 225 357
rect 231 351 237 357
rect 243 351 249 357
rect 255 351 261 357
rect 267 351 273 357
rect 279 351 285 357
rect 291 351 297 357
rect 303 351 309 357
rect 315 351 321 357
rect 327 351 333 357
rect 339 351 345 357
rect 351 351 357 357
rect 363 351 369 357
rect 375 351 381 357
rect 387 351 393 357
rect 399 351 405 357
rect 411 351 417 357
rect 423 351 429 357
rect 435 351 441 357
rect 447 351 453 357
rect 459 351 465 357
rect 471 351 477 357
rect 483 351 489 357
rect 495 351 501 357
rect 507 351 513 357
rect 519 351 525 357
rect 531 351 537 357
rect 543 351 549 357
rect 555 351 561 357
rect 567 351 573 357
rect 579 351 585 357
rect 591 351 597 357
rect 603 351 609 357
rect 615 351 621 357
rect 627 351 633 357
rect 639 351 645 357
rect 651 351 657 357
rect 663 351 669 357
rect 675 351 681 357
rect 687 351 693 357
rect 699 351 705 357
rect 711 351 717 357
rect 723 351 729 357
rect 735 351 741 357
rect 747 351 753 357
rect 759 351 765 357
rect 771 351 777 357
rect 783 351 789 357
rect 795 351 801 357
rect 807 351 813 357
rect 819 351 825 357
rect 831 351 837 357
rect 843 351 849 357
rect 855 351 861 357
rect 867 351 873 357
rect 879 351 885 357
rect 891 351 897 357
rect 903 351 909 357
rect 915 351 921 357
rect 927 351 933 357
rect 939 351 945 357
rect 951 351 957 357
rect 963 351 969 357
rect 975 351 981 357
rect 987 351 993 357
rect 999 351 1005 357
rect 1011 351 1017 357
rect 1023 351 1029 357
rect 1035 351 1041 357
rect 1047 351 1053 357
rect 1059 351 1065 357
rect 1071 351 1077 357
rect 1083 351 1089 357
rect 1095 351 1101 357
rect 1107 351 1113 357
rect 1119 351 1125 357
rect 1131 351 1137 357
rect 1143 351 1149 357
rect 1155 351 1161 357
rect 1167 351 1173 357
rect 1179 351 1185 357
rect 1191 351 1197 357
rect 1203 351 1209 357
rect 1215 351 1221 357
rect 1227 351 1233 357
rect 1239 351 1245 357
rect 1251 351 1257 357
rect 1263 351 1269 357
rect 1275 351 1281 357
rect 1287 351 1293 357
rect 1299 351 1305 357
rect 1311 351 1317 357
rect 1323 351 1329 357
rect 1335 351 1341 357
rect 1347 351 1353 357
rect 1359 351 1365 357
rect 1371 351 1377 357
rect 1383 351 1389 357
rect 1395 351 1401 357
rect 1407 351 1413 357
rect 1419 351 1425 357
rect 1431 351 1437 357
rect 1443 351 1449 357
rect 1455 351 1461 357
rect 1467 351 1473 357
rect 1479 351 1485 357
rect 1491 351 1497 357
rect 1503 351 1509 357
rect 1515 351 1521 357
rect 1527 351 1533 357
rect 1539 351 1545 357
rect 1551 351 1557 357
rect 1563 351 1569 357
rect 1575 351 1581 357
rect 1587 351 1593 357
rect 1599 351 1605 357
<< mvnsubdiffcont >>
rect -57 495 -51 501
rect -45 495 -39 501
rect -33 495 -27 501
rect -21 495 -15 501
rect -9 495 -3 501
rect 3 495 9 501
rect 15 495 21 501
rect 27 495 33 501
rect 39 495 45 501
rect 51 495 57 501
rect 63 495 69 501
rect 75 495 81 501
rect 87 495 93 501
rect 99 495 105 501
rect 111 495 117 501
rect 123 495 129 501
rect 135 495 141 501
rect 147 495 153 501
rect 159 495 165 501
rect 171 495 177 501
rect 183 495 189 501
rect 195 495 201 501
rect 207 495 213 501
rect 219 495 225 501
rect 231 495 237 501
rect 243 495 249 501
rect 255 495 261 501
rect 267 495 273 501
rect 279 495 285 501
rect 291 495 297 501
rect 303 495 309 501
rect 315 495 321 501
rect 327 495 333 501
rect 339 495 345 501
rect 351 495 357 501
rect 363 495 369 501
rect 375 495 381 501
rect 387 495 393 501
rect 399 495 405 501
rect 411 495 417 501
rect 423 495 429 501
rect 435 495 441 501
rect 447 495 453 501
rect 459 495 465 501
rect 471 495 477 501
rect 483 495 489 501
rect 495 495 501 501
rect 507 495 513 501
rect 519 495 525 501
rect 531 495 537 501
rect 543 495 549 501
rect 555 495 561 501
rect 567 495 573 501
rect 579 495 585 501
rect 591 495 597 501
rect 603 495 609 501
rect 615 495 621 501
rect 627 495 633 501
rect 639 495 645 501
rect 651 495 657 501
rect 663 495 669 501
rect 675 495 681 501
rect 687 495 693 501
rect 699 495 705 501
rect 711 495 717 501
rect 723 495 729 501
rect 735 495 741 501
rect 747 495 753 501
rect 759 495 765 501
rect 771 495 777 501
rect 783 495 789 501
rect 795 495 801 501
rect 807 495 813 501
rect 819 495 825 501
rect 831 495 837 501
rect 843 495 849 501
rect 855 495 861 501
rect 867 495 873 501
rect 879 495 885 501
rect 891 495 897 501
rect 903 495 909 501
rect 915 495 921 501
rect 927 495 933 501
rect 939 495 945 501
rect 951 495 957 501
rect 963 495 969 501
rect 975 495 981 501
rect 987 495 993 501
rect 999 495 1005 501
rect 1011 495 1017 501
rect 1023 495 1029 501
rect 1035 495 1041 501
rect 1047 495 1053 501
rect 1059 495 1065 501
rect 1071 495 1077 501
rect 1083 495 1089 501
rect 1095 495 1101 501
rect 1107 495 1113 501
rect 1119 495 1125 501
rect 1131 495 1137 501
rect 1143 495 1149 501
rect 1155 495 1161 501
rect 1167 495 1173 501
rect 1179 495 1185 501
rect 1191 495 1197 501
rect 1203 495 1209 501
rect 1215 495 1221 501
rect 1227 495 1233 501
rect 1239 495 1245 501
rect 1251 495 1257 501
rect 1263 495 1269 501
rect 1275 495 1281 501
rect 1287 495 1293 501
rect 1299 495 1305 501
rect 1311 495 1317 501
rect 1323 495 1329 501
rect 1335 495 1341 501
rect 1347 495 1353 501
rect 1359 495 1365 501
rect 1371 495 1377 501
rect 1383 495 1389 501
rect 1395 495 1401 501
rect 1407 495 1413 501
rect 1419 495 1425 501
rect 1431 495 1437 501
rect 1443 495 1449 501
rect 1455 495 1461 501
rect 1467 495 1473 501
rect 1479 495 1485 501
rect 1491 495 1497 501
rect 1503 495 1509 501
rect 1515 495 1521 501
rect 1527 495 1533 501
rect 1539 495 1545 501
rect 1551 495 1557 501
rect 1563 495 1569 501
rect 1575 495 1581 501
<< polysilicon >>
rect -48 573 -12 576
rect -48 567 -45 573
rect -39 567 -33 573
rect -27 567 -21 573
rect -15 567 -12 573
rect -48 564 -12 567
rect -48 552 -36 564
rect -24 552 -12 564
rect 0 573 36 576
rect 0 567 3 573
rect 9 567 15 573
rect 21 567 27 573
rect 33 567 36 573
rect 0 564 36 567
rect 0 552 12 564
rect 24 552 36 564
rect 48 573 84 576
rect 48 567 51 573
rect 57 567 63 573
rect 69 567 75 573
rect 81 567 84 573
rect 48 564 84 567
rect 48 552 60 564
rect 72 552 84 564
rect 96 573 132 576
rect 96 567 99 573
rect 105 567 111 573
rect 117 567 123 573
rect 129 567 132 573
rect 96 564 132 567
rect 96 552 108 564
rect 120 552 132 564
rect 144 573 180 576
rect 144 567 147 573
rect 153 567 159 573
rect 165 567 171 573
rect 177 567 180 573
rect 144 564 180 567
rect 144 552 156 564
rect 168 552 180 564
rect 192 573 228 576
rect 192 567 195 573
rect 201 567 207 573
rect 213 567 219 573
rect 225 567 228 573
rect 192 564 228 567
rect 192 552 204 564
rect 216 552 228 564
rect 240 573 276 576
rect 240 567 243 573
rect 249 567 255 573
rect 261 567 267 573
rect 273 567 276 573
rect 240 564 276 567
rect 240 552 252 564
rect 264 552 276 564
rect 288 573 324 576
rect 288 567 291 573
rect 297 567 303 573
rect 309 567 315 573
rect 321 567 324 573
rect 288 564 324 567
rect 288 552 300 564
rect 312 552 324 564
rect 336 573 372 576
rect 336 567 339 573
rect 345 567 351 573
rect 357 567 363 573
rect 369 567 372 573
rect 336 564 372 567
rect 336 552 348 564
rect 360 552 372 564
rect 384 573 420 576
rect 384 567 387 573
rect 393 567 399 573
rect 405 567 411 573
rect 417 567 420 573
rect 384 564 420 567
rect 384 552 396 564
rect 408 552 420 564
rect 432 573 468 576
rect 432 567 435 573
rect 441 567 447 573
rect 453 567 459 573
rect 465 567 468 573
rect 432 564 468 567
rect 432 552 444 564
rect 456 552 468 564
rect 480 573 516 576
rect 480 567 483 573
rect 489 567 495 573
rect 501 567 507 573
rect 513 567 516 573
rect 480 564 516 567
rect 480 552 492 564
rect 504 552 516 564
rect 528 573 564 576
rect 528 567 531 573
rect 537 567 543 573
rect 549 567 555 573
rect 561 567 564 573
rect 528 564 564 567
rect 528 552 540 564
rect 552 552 564 564
rect 576 573 612 576
rect 576 567 579 573
rect 585 567 591 573
rect 597 567 603 573
rect 609 567 612 573
rect 576 564 612 567
rect 576 552 588 564
rect 600 552 612 564
rect 624 573 660 576
rect 624 567 627 573
rect 633 567 639 573
rect 645 567 651 573
rect 657 567 660 573
rect 624 564 660 567
rect 624 552 636 564
rect 648 552 660 564
rect 672 573 708 576
rect 672 567 675 573
rect 681 567 687 573
rect 693 567 699 573
rect 705 567 708 573
rect 672 564 708 567
rect 672 552 684 564
rect 696 552 708 564
rect 720 573 756 576
rect 720 567 723 573
rect 729 567 735 573
rect 741 567 747 573
rect 753 567 756 573
rect 720 564 756 567
rect 720 552 732 564
rect 744 552 756 564
rect 768 573 804 576
rect 768 567 771 573
rect 777 567 783 573
rect 789 567 795 573
rect 801 567 804 573
rect 768 564 804 567
rect 768 552 780 564
rect 792 552 804 564
rect 816 573 852 576
rect 816 567 819 573
rect 825 567 831 573
rect 837 567 843 573
rect 849 567 852 573
rect 816 564 852 567
rect 816 552 828 564
rect 840 552 852 564
rect 864 573 900 576
rect 864 567 867 573
rect 873 567 879 573
rect 885 567 891 573
rect 897 567 900 573
rect 864 564 900 567
rect 864 552 876 564
rect 888 552 900 564
rect 912 573 948 576
rect 912 567 915 573
rect 921 567 927 573
rect 933 567 939 573
rect 945 567 948 573
rect 912 564 948 567
rect 912 552 924 564
rect 936 552 948 564
rect 960 573 996 576
rect 960 567 963 573
rect 969 567 975 573
rect 981 567 987 573
rect 993 567 996 573
rect 960 564 996 567
rect 960 552 972 564
rect 984 552 996 564
rect 1008 573 1044 576
rect 1008 567 1011 573
rect 1017 567 1023 573
rect 1029 567 1035 573
rect 1041 567 1044 573
rect 1008 564 1044 567
rect 1008 552 1020 564
rect 1032 552 1044 564
rect 1056 573 1092 576
rect 1056 567 1059 573
rect 1065 567 1071 573
rect 1077 567 1083 573
rect 1089 567 1092 573
rect 1056 564 1092 567
rect 1056 552 1068 564
rect 1080 552 1092 564
rect 1104 573 1140 576
rect 1104 567 1107 573
rect 1113 567 1119 573
rect 1125 567 1131 573
rect 1137 567 1140 573
rect 1104 564 1140 567
rect 1104 552 1116 564
rect 1128 552 1140 564
rect 1152 573 1188 576
rect 1152 567 1155 573
rect 1161 567 1167 573
rect 1173 567 1179 573
rect 1185 567 1188 573
rect 1152 564 1188 567
rect 1152 552 1164 564
rect 1176 552 1188 564
rect 1200 573 1236 576
rect 1200 567 1203 573
rect 1209 567 1215 573
rect 1221 567 1227 573
rect 1233 567 1236 573
rect 1200 564 1236 567
rect 1200 552 1212 564
rect 1224 552 1236 564
rect 1248 573 1284 576
rect 1248 567 1251 573
rect 1257 567 1263 573
rect 1269 567 1275 573
rect 1281 567 1284 573
rect 1248 564 1284 567
rect 1248 552 1260 564
rect 1272 552 1284 564
rect 1296 573 1332 576
rect 1296 567 1299 573
rect 1305 567 1311 573
rect 1317 567 1323 573
rect 1329 567 1332 573
rect 1296 564 1332 567
rect 1296 552 1308 564
rect 1320 552 1332 564
rect 1344 573 1380 576
rect 1344 567 1347 573
rect 1353 567 1359 573
rect 1365 567 1371 573
rect 1377 567 1380 573
rect 1344 564 1380 567
rect 1344 552 1356 564
rect 1368 552 1380 564
rect 1392 573 1428 576
rect 1392 567 1395 573
rect 1401 567 1407 573
rect 1413 567 1419 573
rect 1425 567 1428 573
rect 1392 564 1428 567
rect 1392 552 1404 564
rect 1416 552 1428 564
rect 1440 573 1476 576
rect 1440 567 1443 573
rect 1449 567 1455 573
rect 1461 567 1467 573
rect 1473 567 1476 573
rect 1440 564 1476 567
rect 1440 552 1452 564
rect 1464 552 1476 564
rect 1488 573 1524 576
rect 1488 567 1491 573
rect 1497 567 1503 573
rect 1509 567 1515 573
rect 1521 567 1524 573
rect 1488 564 1524 567
rect 1488 552 1500 564
rect 1512 552 1524 564
rect 1536 573 1572 576
rect 1536 567 1539 573
rect 1545 567 1551 573
rect 1557 567 1563 573
rect 1569 567 1572 573
rect 1536 564 1572 567
rect 1536 552 1548 564
rect 1560 552 1572 564
rect -48 510 -36 516
rect -24 510 -12 516
rect 0 510 12 516
rect 24 510 36 516
rect 48 510 60 516
rect 72 510 84 516
rect 96 510 108 516
rect 120 510 132 516
rect 144 510 156 516
rect 168 510 180 516
rect 192 510 204 516
rect 216 510 228 516
rect 240 510 252 516
rect 264 510 276 516
rect 288 510 300 516
rect 312 510 324 516
rect 336 510 348 516
rect 360 510 372 516
rect 384 510 396 516
rect 408 510 420 516
rect 432 510 444 516
rect 456 510 468 516
rect 480 510 492 516
rect 504 510 516 516
rect 528 510 540 516
rect 552 510 564 516
rect 576 510 588 516
rect 600 510 612 516
rect 624 510 636 516
rect 648 510 660 516
rect 672 510 684 516
rect 696 510 708 516
rect 720 510 732 516
rect 744 510 756 516
rect 768 510 780 516
rect 792 510 804 516
rect 816 510 828 516
rect 840 510 852 516
rect 864 510 876 516
rect 888 510 900 516
rect 912 510 924 516
rect 936 510 948 516
rect 960 510 972 516
rect 984 510 996 516
rect 1008 510 1020 516
rect 1032 510 1044 516
rect 1056 510 1068 516
rect 1080 510 1092 516
rect 1104 510 1116 516
rect 1128 510 1140 516
rect 1152 510 1164 516
rect 1176 510 1188 516
rect 1200 510 1212 516
rect 1224 510 1236 516
rect 1248 510 1260 516
rect 1272 510 1284 516
rect 1296 510 1308 516
rect 1320 510 1332 516
rect 1344 510 1356 516
rect 1368 510 1380 516
rect 1392 510 1404 516
rect 1416 510 1428 516
rect 1440 510 1452 516
rect 1464 510 1476 516
rect 1488 510 1500 516
rect 1512 510 1524 516
rect 1536 510 1548 516
rect 1560 510 1572 516
rect -48 426 -36 432
rect -24 426 -12 432
rect 0 426 12 432
rect 24 426 36 432
rect 48 426 60 432
rect 72 426 84 432
rect 96 426 108 432
rect 120 426 132 432
rect 144 426 156 432
rect 168 426 180 432
rect 192 426 204 432
rect 216 426 228 432
rect 240 426 252 432
rect 264 426 276 432
rect 288 426 300 432
rect 312 426 324 432
rect 336 426 348 432
rect 360 426 372 432
rect 384 426 396 432
rect 408 426 420 432
rect 432 426 444 432
rect 456 426 468 432
rect 480 426 492 432
rect 504 426 516 432
rect 528 426 540 432
rect 552 426 564 432
rect 576 426 588 432
rect 600 426 612 432
rect 624 426 636 432
rect 648 426 660 432
rect 672 426 684 432
rect 696 426 708 432
rect 720 426 732 432
rect 744 426 756 432
rect 768 426 780 432
rect 792 426 804 432
rect 816 426 828 432
rect 840 426 852 432
rect 864 426 876 432
rect 888 426 900 432
rect 912 426 924 432
rect 936 426 948 432
rect 960 426 972 432
rect 984 426 996 432
rect 1008 426 1020 432
rect 1032 426 1044 432
rect 1056 426 1068 432
rect 1080 426 1092 432
rect 1104 426 1116 432
rect 1128 426 1140 432
rect 1152 426 1164 432
rect 1176 426 1188 432
rect 1200 426 1212 432
rect 1224 426 1236 432
rect 1248 426 1260 432
rect 1272 426 1284 432
rect 1296 426 1308 432
rect 1320 426 1332 432
rect 1344 426 1356 432
rect 1368 426 1380 432
rect 1392 426 1404 432
rect 1416 426 1428 432
rect 1440 426 1452 432
rect 1464 426 1476 432
rect 1488 426 1500 432
rect 1512 426 1524 432
rect 1536 426 1548 432
rect 1560 426 1572 432
rect -48 384 -36 396
rect -24 384 -12 396
rect -48 381 -12 384
rect -48 375 -45 381
rect -39 375 -33 381
rect -27 375 -21 381
rect -15 375 -12 381
rect -48 372 -12 375
rect 0 384 12 396
rect 24 384 36 396
rect 0 381 36 384
rect 0 375 3 381
rect 9 375 15 381
rect 21 375 27 381
rect 33 375 36 381
rect 0 372 36 375
rect 48 384 60 396
rect 72 384 84 396
rect 48 381 84 384
rect 48 375 51 381
rect 57 375 63 381
rect 69 375 75 381
rect 81 375 84 381
rect 48 372 84 375
rect 96 384 108 396
rect 120 384 132 396
rect 96 381 132 384
rect 96 375 99 381
rect 105 375 111 381
rect 117 375 123 381
rect 129 375 132 381
rect 96 372 132 375
rect 144 384 156 396
rect 168 384 180 396
rect 144 381 180 384
rect 144 375 147 381
rect 153 375 159 381
rect 165 375 171 381
rect 177 375 180 381
rect 144 372 180 375
rect 192 384 204 396
rect 216 384 228 396
rect 192 381 228 384
rect 192 375 195 381
rect 201 375 207 381
rect 213 375 219 381
rect 225 375 228 381
rect 192 372 228 375
rect 240 384 252 396
rect 264 384 276 396
rect 240 381 276 384
rect 240 375 243 381
rect 249 375 255 381
rect 261 375 267 381
rect 273 375 276 381
rect 240 372 276 375
rect 288 384 300 396
rect 312 384 324 396
rect 288 381 324 384
rect 288 375 291 381
rect 297 375 303 381
rect 309 375 315 381
rect 321 375 324 381
rect 288 372 324 375
rect 336 384 348 396
rect 360 384 372 396
rect 336 381 372 384
rect 336 375 339 381
rect 345 375 351 381
rect 357 375 363 381
rect 369 375 372 381
rect 336 372 372 375
rect 384 384 396 396
rect 408 384 420 396
rect 384 381 420 384
rect 384 375 387 381
rect 393 375 399 381
rect 405 375 411 381
rect 417 375 420 381
rect 384 372 420 375
rect 432 384 444 396
rect 456 384 468 396
rect 432 381 468 384
rect 432 375 435 381
rect 441 375 447 381
rect 453 375 459 381
rect 465 375 468 381
rect 432 372 468 375
rect 480 384 492 396
rect 504 384 516 396
rect 480 381 516 384
rect 480 375 483 381
rect 489 375 495 381
rect 501 375 507 381
rect 513 375 516 381
rect 480 372 516 375
rect 528 384 540 396
rect 552 384 564 396
rect 528 381 564 384
rect 528 375 531 381
rect 537 375 543 381
rect 549 375 555 381
rect 561 375 564 381
rect 528 372 564 375
rect 576 384 588 396
rect 600 384 612 396
rect 576 381 612 384
rect 576 375 579 381
rect 585 375 591 381
rect 597 375 603 381
rect 609 375 612 381
rect 576 372 612 375
rect 624 384 636 396
rect 648 384 660 396
rect 624 381 660 384
rect 624 375 627 381
rect 633 375 639 381
rect 645 375 651 381
rect 657 375 660 381
rect 624 372 660 375
rect 672 384 684 396
rect 696 384 708 396
rect 672 381 708 384
rect 672 375 675 381
rect 681 375 687 381
rect 693 375 699 381
rect 705 375 708 381
rect 672 372 708 375
rect 720 384 732 396
rect 744 384 756 396
rect 720 381 756 384
rect 720 375 723 381
rect 729 375 735 381
rect 741 375 747 381
rect 753 375 756 381
rect 720 372 756 375
rect 768 384 780 396
rect 792 384 804 396
rect 768 381 804 384
rect 768 375 771 381
rect 777 375 783 381
rect 789 375 795 381
rect 801 375 804 381
rect 768 372 804 375
rect 816 384 828 396
rect 840 384 852 396
rect 816 381 852 384
rect 816 375 819 381
rect 825 375 831 381
rect 837 375 843 381
rect 849 375 852 381
rect 816 372 852 375
rect 864 384 876 396
rect 888 384 900 396
rect 864 381 900 384
rect 864 375 867 381
rect 873 375 879 381
rect 885 375 891 381
rect 897 375 900 381
rect 864 372 900 375
rect 912 384 924 396
rect 936 384 948 396
rect 912 381 948 384
rect 912 375 915 381
rect 921 375 927 381
rect 933 375 939 381
rect 945 375 948 381
rect 912 372 948 375
rect 960 384 972 396
rect 984 384 996 396
rect 960 381 996 384
rect 960 375 963 381
rect 969 375 975 381
rect 981 375 987 381
rect 993 375 996 381
rect 960 372 996 375
rect 1008 384 1020 396
rect 1032 384 1044 396
rect 1008 381 1044 384
rect 1008 375 1011 381
rect 1017 375 1023 381
rect 1029 375 1035 381
rect 1041 375 1044 381
rect 1008 372 1044 375
rect 1056 384 1068 396
rect 1080 384 1092 396
rect 1056 381 1092 384
rect 1056 375 1059 381
rect 1065 375 1071 381
rect 1077 375 1083 381
rect 1089 375 1092 381
rect 1056 372 1092 375
rect 1104 384 1116 396
rect 1128 384 1140 396
rect 1104 381 1140 384
rect 1104 375 1107 381
rect 1113 375 1119 381
rect 1125 375 1131 381
rect 1137 375 1140 381
rect 1104 372 1140 375
rect 1152 384 1164 396
rect 1176 384 1188 396
rect 1152 381 1188 384
rect 1152 375 1155 381
rect 1161 375 1167 381
rect 1173 375 1179 381
rect 1185 375 1188 381
rect 1152 372 1188 375
rect 1200 384 1212 396
rect 1224 384 1236 396
rect 1200 381 1236 384
rect 1200 375 1203 381
rect 1209 375 1215 381
rect 1221 375 1227 381
rect 1233 375 1236 381
rect 1200 372 1236 375
rect 1248 384 1260 396
rect 1272 384 1284 396
rect 1248 381 1284 384
rect 1248 375 1251 381
rect 1257 375 1263 381
rect 1269 375 1275 381
rect 1281 375 1284 381
rect 1248 372 1284 375
rect 1296 384 1308 396
rect 1320 384 1332 396
rect 1296 381 1332 384
rect 1296 375 1299 381
rect 1305 375 1311 381
rect 1317 375 1323 381
rect 1329 375 1332 381
rect 1296 372 1332 375
rect 1344 384 1356 396
rect 1368 384 1380 396
rect 1344 381 1380 384
rect 1344 375 1347 381
rect 1353 375 1359 381
rect 1365 375 1371 381
rect 1377 375 1380 381
rect 1344 372 1380 375
rect 1392 384 1404 396
rect 1416 384 1428 396
rect 1392 381 1428 384
rect 1392 375 1395 381
rect 1401 375 1407 381
rect 1413 375 1419 381
rect 1425 375 1428 381
rect 1392 372 1428 375
rect 1440 384 1452 396
rect 1464 384 1476 396
rect 1440 381 1476 384
rect 1440 375 1443 381
rect 1449 375 1455 381
rect 1461 375 1467 381
rect 1473 375 1476 381
rect 1440 372 1476 375
rect 1488 384 1500 396
rect 1512 384 1524 396
rect 1488 381 1524 384
rect 1488 375 1491 381
rect 1497 375 1503 381
rect 1509 375 1515 381
rect 1521 375 1524 381
rect 1488 372 1524 375
rect 1536 384 1548 396
rect 1560 384 1572 396
rect 1536 381 1572 384
rect 1536 375 1539 381
rect 1545 375 1551 381
rect 1557 375 1563 381
rect 1569 375 1572 381
rect 1536 372 1572 375
rect -48 69 -12 72
rect -48 63 -45 69
rect -39 63 -33 69
rect -27 63 -21 69
rect -15 63 -12 69
rect -48 60 -12 63
rect -48 48 -36 60
rect -24 48 -12 60
rect 0 69 36 72
rect 0 63 3 69
rect 9 63 15 69
rect 21 63 27 69
rect 33 63 36 69
rect 0 60 36 63
rect 0 48 12 60
rect 24 48 36 60
rect 48 69 84 72
rect 48 63 51 69
rect 57 63 63 69
rect 69 63 75 69
rect 81 63 84 69
rect 48 60 84 63
rect 48 48 60 60
rect 72 48 84 60
rect 96 69 132 72
rect 96 63 99 69
rect 105 63 111 69
rect 117 63 123 69
rect 129 63 132 69
rect 96 60 132 63
rect 96 48 108 60
rect 120 48 132 60
rect 144 69 180 72
rect 144 63 147 69
rect 153 63 159 69
rect 165 63 171 69
rect 177 63 180 69
rect 144 60 180 63
rect 144 48 156 60
rect 168 48 180 60
rect 192 69 228 72
rect 192 63 195 69
rect 201 63 207 69
rect 213 63 219 69
rect 225 63 228 69
rect 192 60 228 63
rect 192 48 204 60
rect 216 48 228 60
rect 240 69 276 72
rect 240 63 243 69
rect 249 63 255 69
rect 261 63 267 69
rect 273 63 276 69
rect 240 60 276 63
rect 240 48 252 60
rect 264 48 276 60
rect 288 69 324 72
rect 288 63 291 69
rect 297 63 303 69
rect 309 63 315 69
rect 321 63 324 69
rect 288 60 324 63
rect 288 48 300 60
rect 312 48 324 60
rect 336 69 372 72
rect 336 63 339 69
rect 345 63 351 69
rect 357 63 363 69
rect 369 63 372 69
rect 336 60 372 63
rect 336 48 348 60
rect 360 48 372 60
rect 384 69 420 72
rect 384 63 387 69
rect 393 63 399 69
rect 405 63 411 69
rect 417 63 420 69
rect 384 60 420 63
rect 384 48 396 60
rect 408 48 420 60
rect 432 69 468 72
rect 432 63 435 69
rect 441 63 447 69
rect 453 63 459 69
rect 465 63 468 69
rect 432 60 468 63
rect 432 48 444 60
rect 456 48 468 60
rect 480 69 516 72
rect 480 63 483 69
rect 489 63 495 69
rect 501 63 507 69
rect 513 63 516 69
rect 480 60 516 63
rect 480 48 492 60
rect 504 48 516 60
rect 528 69 564 72
rect 528 63 531 69
rect 537 63 543 69
rect 549 63 555 69
rect 561 63 564 69
rect 528 60 564 63
rect 528 48 540 60
rect 552 48 564 60
rect 576 69 612 72
rect 576 63 579 69
rect 585 63 591 69
rect 597 63 603 69
rect 609 63 612 69
rect 576 60 612 63
rect 576 48 588 60
rect 600 48 612 60
rect 624 69 660 72
rect 624 63 627 69
rect 633 63 639 69
rect 645 63 651 69
rect 657 63 660 69
rect 624 60 660 63
rect 624 48 636 60
rect 648 48 660 60
rect 672 69 708 72
rect 672 63 675 69
rect 681 63 687 69
rect 693 63 699 69
rect 705 63 708 69
rect 672 60 708 63
rect 672 48 684 60
rect 696 48 708 60
rect 720 69 756 72
rect 720 63 723 69
rect 729 63 735 69
rect 741 63 747 69
rect 753 63 756 69
rect 720 60 756 63
rect 720 48 732 60
rect 744 48 756 60
rect 768 69 804 72
rect 768 63 771 69
rect 777 63 783 69
rect 789 63 795 69
rect 801 63 804 69
rect 768 60 804 63
rect 768 48 780 60
rect 792 48 804 60
rect 816 69 852 72
rect 816 63 819 69
rect 825 63 831 69
rect 837 63 843 69
rect 849 63 852 69
rect 816 60 852 63
rect 816 48 828 60
rect 840 48 852 60
rect 864 69 900 72
rect 864 63 867 69
rect 873 63 879 69
rect 885 63 891 69
rect 897 63 900 69
rect 864 60 900 63
rect 864 48 876 60
rect 888 48 900 60
rect 912 69 948 72
rect 912 63 915 69
rect 921 63 927 69
rect 933 63 939 69
rect 945 63 948 69
rect 912 60 948 63
rect 912 48 924 60
rect 936 48 948 60
rect 960 69 996 72
rect 960 63 963 69
rect 969 63 975 69
rect 981 63 987 69
rect 993 63 996 69
rect 960 60 996 63
rect 960 48 972 60
rect 984 48 996 60
rect 1008 69 1044 72
rect 1008 63 1011 69
rect 1017 63 1023 69
rect 1029 63 1035 69
rect 1041 63 1044 69
rect 1008 60 1044 63
rect 1008 48 1020 60
rect 1032 48 1044 60
rect 1056 69 1092 72
rect 1056 63 1059 69
rect 1065 63 1071 69
rect 1077 63 1083 69
rect 1089 63 1092 69
rect 1056 60 1092 63
rect 1056 48 1068 60
rect 1080 48 1092 60
rect 1104 69 1140 72
rect 1104 63 1107 69
rect 1113 63 1119 69
rect 1125 63 1131 69
rect 1137 63 1140 69
rect 1104 60 1140 63
rect 1104 48 1116 60
rect 1128 48 1140 60
rect 1152 69 1188 72
rect 1152 63 1155 69
rect 1161 63 1167 69
rect 1173 63 1179 69
rect 1185 63 1188 69
rect 1152 60 1188 63
rect 1152 48 1164 60
rect 1176 48 1188 60
rect 1200 69 1236 72
rect 1200 63 1203 69
rect 1209 63 1215 69
rect 1221 63 1227 69
rect 1233 63 1236 69
rect 1200 60 1236 63
rect 1200 48 1212 60
rect 1224 48 1236 60
rect 1248 69 1284 72
rect 1248 63 1251 69
rect 1257 63 1263 69
rect 1269 63 1275 69
rect 1281 63 1284 69
rect 1248 60 1284 63
rect 1248 48 1260 60
rect 1272 48 1284 60
rect 1296 69 1332 72
rect 1296 63 1299 69
rect 1305 63 1311 69
rect 1317 63 1323 69
rect 1329 63 1332 69
rect 1296 60 1332 63
rect 1296 48 1308 60
rect 1320 48 1332 60
rect 1344 69 1380 72
rect 1344 63 1347 69
rect 1353 63 1359 69
rect 1365 63 1371 69
rect 1377 63 1380 69
rect 1344 60 1380 63
rect 1344 48 1356 60
rect 1368 48 1380 60
rect 1392 69 1428 72
rect 1392 63 1395 69
rect 1401 63 1407 69
rect 1413 63 1419 69
rect 1425 63 1428 69
rect 1392 60 1428 63
rect 1392 48 1404 60
rect 1416 48 1428 60
rect 1440 69 1476 72
rect 1440 63 1443 69
rect 1449 63 1455 69
rect 1461 63 1467 69
rect 1473 63 1476 69
rect 1440 60 1476 63
rect 1440 48 1452 60
rect 1464 48 1476 60
rect 1488 69 1524 72
rect 1488 63 1491 69
rect 1497 63 1503 69
rect 1509 63 1515 69
rect 1521 63 1524 69
rect 1488 60 1524 63
rect 1488 48 1500 60
rect 1512 48 1524 60
rect 1536 69 1572 72
rect 1536 63 1539 69
rect 1545 63 1551 69
rect 1557 63 1563 69
rect 1569 63 1572 69
rect 1536 60 1572 63
rect 1536 48 1548 60
rect 1560 48 1572 60
rect -48 6 -36 12
rect -24 6 -12 12
rect 0 6 12 12
rect 24 6 36 12
rect 48 6 60 12
rect 72 6 84 12
rect 96 6 108 12
rect 120 6 132 12
rect 144 6 156 12
rect 168 6 180 12
rect 192 6 204 12
rect 216 6 228 12
rect 240 6 252 12
rect 264 6 276 12
rect 288 6 300 12
rect 312 6 324 12
rect 336 6 348 12
rect 360 6 372 12
rect 384 6 396 12
rect 408 6 420 12
rect 432 6 444 12
rect 456 6 468 12
rect 480 6 492 12
rect 504 6 516 12
rect 528 6 540 12
rect 552 6 564 12
rect 576 6 588 12
rect 600 6 612 12
rect 624 6 636 12
rect 648 6 660 12
rect 672 6 684 12
rect 696 6 708 12
rect 720 6 732 12
rect 744 6 756 12
rect 768 6 780 12
rect 792 6 804 12
rect 816 6 828 12
rect 840 6 852 12
rect 864 6 876 12
rect 888 6 900 12
rect 912 6 924 12
rect 936 6 948 12
rect 960 6 972 12
rect 984 6 996 12
rect 1008 6 1020 12
rect 1032 6 1044 12
rect 1056 6 1068 12
rect 1080 6 1092 12
rect 1104 6 1116 12
rect 1128 6 1140 12
rect 1152 6 1164 12
rect 1176 6 1188 12
rect 1200 6 1212 12
rect 1224 6 1236 12
rect 1248 6 1260 12
rect 1272 6 1284 12
rect 1296 6 1308 12
rect 1320 6 1332 12
rect 1344 6 1356 12
rect 1368 6 1380 12
rect 1392 6 1404 12
rect 1416 6 1428 12
rect 1440 6 1452 12
rect 1464 6 1476 12
rect 1488 6 1500 12
rect 1512 6 1524 12
rect 1536 6 1548 12
rect 1560 6 1572 12
<< polycontact >>
rect -45 567 -39 573
rect -33 567 -27 573
rect -21 567 -15 573
rect 3 567 9 573
rect 15 567 21 573
rect 27 567 33 573
rect 51 567 57 573
rect 63 567 69 573
rect 75 567 81 573
rect 99 567 105 573
rect 111 567 117 573
rect 123 567 129 573
rect 147 567 153 573
rect 159 567 165 573
rect 171 567 177 573
rect 195 567 201 573
rect 207 567 213 573
rect 219 567 225 573
rect 243 567 249 573
rect 255 567 261 573
rect 267 567 273 573
rect 291 567 297 573
rect 303 567 309 573
rect 315 567 321 573
rect 339 567 345 573
rect 351 567 357 573
rect 363 567 369 573
rect 387 567 393 573
rect 399 567 405 573
rect 411 567 417 573
rect 435 567 441 573
rect 447 567 453 573
rect 459 567 465 573
rect 483 567 489 573
rect 495 567 501 573
rect 507 567 513 573
rect 531 567 537 573
rect 543 567 549 573
rect 555 567 561 573
rect 579 567 585 573
rect 591 567 597 573
rect 603 567 609 573
rect 627 567 633 573
rect 639 567 645 573
rect 651 567 657 573
rect 675 567 681 573
rect 687 567 693 573
rect 699 567 705 573
rect 723 567 729 573
rect 735 567 741 573
rect 747 567 753 573
rect 771 567 777 573
rect 783 567 789 573
rect 795 567 801 573
rect 819 567 825 573
rect 831 567 837 573
rect 843 567 849 573
rect 867 567 873 573
rect 879 567 885 573
rect 891 567 897 573
rect 915 567 921 573
rect 927 567 933 573
rect 939 567 945 573
rect 963 567 969 573
rect 975 567 981 573
rect 987 567 993 573
rect 1011 567 1017 573
rect 1023 567 1029 573
rect 1035 567 1041 573
rect 1059 567 1065 573
rect 1071 567 1077 573
rect 1083 567 1089 573
rect 1107 567 1113 573
rect 1119 567 1125 573
rect 1131 567 1137 573
rect 1155 567 1161 573
rect 1167 567 1173 573
rect 1179 567 1185 573
rect 1203 567 1209 573
rect 1215 567 1221 573
rect 1227 567 1233 573
rect 1251 567 1257 573
rect 1263 567 1269 573
rect 1275 567 1281 573
rect 1299 567 1305 573
rect 1311 567 1317 573
rect 1323 567 1329 573
rect 1347 567 1353 573
rect 1359 567 1365 573
rect 1371 567 1377 573
rect 1395 567 1401 573
rect 1407 567 1413 573
rect 1419 567 1425 573
rect 1443 567 1449 573
rect 1455 567 1461 573
rect 1467 567 1473 573
rect 1491 567 1497 573
rect 1503 567 1509 573
rect 1515 567 1521 573
rect 1539 567 1545 573
rect 1551 567 1557 573
rect 1563 567 1569 573
rect -45 375 -39 381
rect -33 375 -27 381
rect -21 375 -15 381
rect 3 375 9 381
rect 15 375 21 381
rect 27 375 33 381
rect 51 375 57 381
rect 63 375 69 381
rect 75 375 81 381
rect 99 375 105 381
rect 111 375 117 381
rect 123 375 129 381
rect 147 375 153 381
rect 159 375 165 381
rect 171 375 177 381
rect 195 375 201 381
rect 207 375 213 381
rect 219 375 225 381
rect 243 375 249 381
rect 255 375 261 381
rect 267 375 273 381
rect 291 375 297 381
rect 303 375 309 381
rect 315 375 321 381
rect 339 375 345 381
rect 351 375 357 381
rect 363 375 369 381
rect 387 375 393 381
rect 399 375 405 381
rect 411 375 417 381
rect 435 375 441 381
rect 447 375 453 381
rect 459 375 465 381
rect 483 375 489 381
rect 495 375 501 381
rect 507 375 513 381
rect 531 375 537 381
rect 543 375 549 381
rect 555 375 561 381
rect 579 375 585 381
rect 591 375 597 381
rect 603 375 609 381
rect 627 375 633 381
rect 639 375 645 381
rect 651 375 657 381
rect 675 375 681 381
rect 687 375 693 381
rect 699 375 705 381
rect 723 375 729 381
rect 735 375 741 381
rect 747 375 753 381
rect 771 375 777 381
rect 783 375 789 381
rect 795 375 801 381
rect 819 375 825 381
rect 831 375 837 381
rect 843 375 849 381
rect 867 375 873 381
rect 879 375 885 381
rect 891 375 897 381
rect 915 375 921 381
rect 927 375 933 381
rect 939 375 945 381
rect 963 375 969 381
rect 975 375 981 381
rect 987 375 993 381
rect 1011 375 1017 381
rect 1023 375 1029 381
rect 1035 375 1041 381
rect 1059 375 1065 381
rect 1071 375 1077 381
rect 1083 375 1089 381
rect 1107 375 1113 381
rect 1119 375 1125 381
rect 1131 375 1137 381
rect 1155 375 1161 381
rect 1167 375 1173 381
rect 1179 375 1185 381
rect 1203 375 1209 381
rect 1215 375 1221 381
rect 1227 375 1233 381
rect 1251 375 1257 381
rect 1263 375 1269 381
rect 1275 375 1281 381
rect 1299 375 1305 381
rect 1311 375 1317 381
rect 1323 375 1329 381
rect 1347 375 1353 381
rect 1359 375 1365 381
rect 1371 375 1377 381
rect 1395 375 1401 381
rect 1407 375 1413 381
rect 1419 375 1425 381
rect 1443 375 1449 381
rect 1455 375 1461 381
rect 1467 375 1473 381
rect 1491 375 1497 381
rect 1503 375 1509 381
rect 1515 375 1521 381
rect 1539 375 1545 381
rect 1551 375 1557 381
rect 1563 375 1569 381
rect -45 63 -39 69
rect -33 63 -27 69
rect -21 63 -15 69
rect 3 63 9 69
rect 15 63 21 69
rect 27 63 33 69
rect 51 63 57 69
rect 63 63 69 69
rect 75 63 81 69
rect 99 63 105 69
rect 111 63 117 69
rect 123 63 129 69
rect 147 63 153 69
rect 159 63 165 69
rect 171 63 177 69
rect 195 63 201 69
rect 207 63 213 69
rect 219 63 225 69
rect 243 63 249 69
rect 255 63 261 69
rect 267 63 273 69
rect 291 63 297 69
rect 303 63 309 69
rect 315 63 321 69
rect 339 63 345 69
rect 351 63 357 69
rect 363 63 369 69
rect 387 63 393 69
rect 399 63 405 69
rect 411 63 417 69
rect 435 63 441 69
rect 447 63 453 69
rect 459 63 465 69
rect 483 63 489 69
rect 495 63 501 69
rect 507 63 513 69
rect 531 63 537 69
rect 543 63 549 69
rect 555 63 561 69
rect 579 63 585 69
rect 591 63 597 69
rect 603 63 609 69
rect 627 63 633 69
rect 639 63 645 69
rect 651 63 657 69
rect 675 63 681 69
rect 687 63 693 69
rect 699 63 705 69
rect 723 63 729 69
rect 735 63 741 69
rect 747 63 753 69
rect 771 63 777 69
rect 783 63 789 69
rect 795 63 801 69
rect 819 63 825 69
rect 831 63 837 69
rect 843 63 849 69
rect 867 63 873 69
rect 879 63 885 69
rect 891 63 897 69
rect 915 63 921 69
rect 927 63 933 69
rect 939 63 945 69
rect 963 63 969 69
rect 975 63 981 69
rect 987 63 993 69
rect 1011 63 1017 69
rect 1023 63 1029 69
rect 1035 63 1041 69
rect 1059 63 1065 69
rect 1071 63 1077 69
rect 1083 63 1089 69
rect 1107 63 1113 69
rect 1119 63 1125 69
rect 1131 63 1137 69
rect 1155 63 1161 69
rect 1167 63 1173 69
rect 1179 63 1185 69
rect 1203 63 1209 69
rect 1215 63 1221 69
rect 1227 63 1233 69
rect 1251 63 1257 69
rect 1263 63 1269 69
rect 1275 63 1281 69
rect 1299 63 1305 69
rect 1311 63 1317 69
rect 1323 63 1329 69
rect 1347 63 1353 69
rect 1359 63 1365 69
rect 1371 63 1377 69
rect 1395 63 1401 69
rect 1407 63 1413 69
rect 1419 63 1425 69
rect 1443 63 1449 69
rect 1455 63 1461 69
rect 1467 63 1473 69
rect 1491 63 1497 69
rect 1503 63 1509 69
rect 1515 63 1521 69
rect 1539 63 1545 69
rect 1551 63 1557 69
rect 1563 63 1569 69
<< metal1 >>
rect -108 621 1632 624
rect -108 615 -105 621
rect -99 615 -93 621
rect -87 615 -81 621
rect -75 615 -69 621
rect -63 615 -57 621
rect -51 615 -45 621
rect -39 615 -33 621
rect -27 615 -21 621
rect -15 615 -9 621
rect -3 615 3 621
rect 9 615 15 621
rect 21 615 27 621
rect 33 615 39 621
rect 45 615 51 621
rect 57 615 63 621
rect 69 615 75 621
rect 81 615 87 621
rect 93 615 99 621
rect 105 615 111 621
rect 117 615 123 621
rect 129 615 135 621
rect 141 615 147 621
rect 153 615 159 621
rect 165 615 171 621
rect 177 615 183 621
rect 189 615 195 621
rect 201 615 207 621
rect 213 615 219 621
rect 225 615 231 621
rect 237 615 243 621
rect 249 615 255 621
rect 261 615 267 621
rect 273 615 279 621
rect 285 615 291 621
rect 297 615 303 621
rect 309 615 315 621
rect 321 615 327 621
rect 333 615 339 621
rect 345 615 351 621
rect 357 615 363 621
rect 369 615 375 621
rect 381 615 387 621
rect 393 615 399 621
rect 405 615 411 621
rect 417 615 423 621
rect 429 615 435 621
rect 441 615 447 621
rect 453 615 459 621
rect 465 615 471 621
rect 477 615 483 621
rect 489 615 495 621
rect 501 615 507 621
rect 513 615 519 621
rect 525 615 531 621
rect 537 615 543 621
rect 549 615 555 621
rect 561 615 567 621
rect 573 615 579 621
rect 585 615 591 621
rect 597 615 603 621
rect 609 615 615 621
rect 621 615 627 621
rect 633 615 639 621
rect 645 615 651 621
rect 657 615 663 621
rect 669 615 675 621
rect 681 615 687 621
rect 693 615 699 621
rect 705 615 711 621
rect 717 615 723 621
rect 729 615 735 621
rect 741 615 747 621
rect 753 615 759 621
rect 765 615 771 621
rect 777 615 783 621
rect 789 615 795 621
rect 801 615 807 621
rect 813 615 819 621
rect 825 615 831 621
rect 837 615 843 621
rect 849 615 855 621
rect 861 615 867 621
rect 873 615 879 621
rect 885 615 891 621
rect 897 615 903 621
rect 909 615 915 621
rect 921 615 927 621
rect 933 615 939 621
rect 945 615 951 621
rect 957 615 963 621
rect 969 615 975 621
rect 981 615 987 621
rect 993 615 999 621
rect 1005 615 1011 621
rect 1017 615 1023 621
rect 1029 615 1035 621
rect 1041 615 1047 621
rect 1053 615 1059 621
rect 1065 615 1071 621
rect 1077 615 1083 621
rect 1089 615 1095 621
rect 1101 615 1107 621
rect 1113 615 1119 621
rect 1125 615 1131 621
rect 1137 615 1143 621
rect 1149 615 1155 621
rect 1161 615 1167 621
rect 1173 615 1179 621
rect 1185 615 1191 621
rect 1197 615 1203 621
rect 1209 615 1215 621
rect 1221 615 1227 621
rect 1233 615 1239 621
rect 1245 615 1251 621
rect 1257 615 1263 621
rect 1269 615 1275 621
rect 1281 615 1287 621
rect 1293 615 1299 621
rect 1305 615 1311 621
rect 1317 615 1323 621
rect 1329 615 1335 621
rect 1341 615 1347 621
rect 1353 615 1359 621
rect 1365 615 1371 621
rect 1377 615 1383 621
rect 1389 615 1395 621
rect 1401 615 1407 621
rect 1413 615 1419 621
rect 1425 615 1431 621
rect 1437 615 1443 621
rect 1449 615 1455 621
rect 1461 615 1467 621
rect 1473 615 1479 621
rect 1485 615 1491 621
rect 1497 615 1503 621
rect 1509 615 1515 621
rect 1521 615 1527 621
rect 1533 615 1539 621
rect 1545 615 1551 621
rect 1557 615 1563 621
rect 1569 615 1575 621
rect 1581 615 1587 621
rect 1593 615 1599 621
rect 1605 615 1611 621
rect 1617 615 1623 621
rect 1629 615 1632 621
rect -108 612 1632 615
rect -108 609 -96 612
rect -108 603 -105 609
rect -99 603 -96 609
rect -108 597 -96 603
rect 1620 609 1632 612
rect 1620 603 1623 609
rect 1629 603 1632 609
rect -108 591 -105 597
rect -99 591 -96 597
rect -108 585 -96 591
rect -108 579 -105 585
rect -99 579 -96 585
rect -108 573 -96 579
rect -108 567 -105 573
rect -99 567 -96 573
rect -108 561 -96 567
rect -108 555 -105 561
rect -99 555 -96 561
rect -108 549 -96 555
rect -108 543 -105 549
rect -99 543 -96 549
rect -108 537 -96 543
rect -108 531 -105 537
rect -99 531 -96 537
rect -108 525 -96 531
rect -108 519 -105 525
rect -99 519 -96 525
rect -108 513 -96 519
rect -108 507 -105 513
rect -99 507 -96 513
rect -108 501 -96 507
rect -108 495 -105 501
rect -99 495 -96 501
rect -108 489 -96 495
rect -84 597 1608 600
rect -84 591 -81 597
rect -75 591 -69 597
rect -63 591 -57 597
rect -51 591 -45 597
rect -39 591 -33 597
rect -27 591 -21 597
rect -15 591 -9 597
rect -3 591 3 597
rect 9 591 15 597
rect 21 591 27 597
rect 33 591 39 597
rect 45 591 51 597
rect 57 591 63 597
rect 69 591 75 597
rect 81 591 87 597
rect 93 591 99 597
rect 105 591 111 597
rect 117 591 123 597
rect 129 591 135 597
rect 141 591 147 597
rect 153 591 159 597
rect 165 591 171 597
rect 177 591 183 597
rect 189 591 195 597
rect 201 591 207 597
rect 213 591 219 597
rect 225 591 231 597
rect 237 591 243 597
rect 249 591 255 597
rect 261 591 267 597
rect 273 591 279 597
rect 285 591 291 597
rect 297 591 303 597
rect 309 591 315 597
rect 321 591 327 597
rect 333 591 339 597
rect 345 591 351 597
rect 357 591 363 597
rect 369 591 375 597
rect 381 591 387 597
rect 393 591 399 597
rect 405 591 411 597
rect 417 591 423 597
rect 429 591 435 597
rect 441 591 447 597
rect 453 591 459 597
rect 465 591 471 597
rect 477 591 483 597
rect 489 591 495 597
rect 501 591 507 597
rect 513 591 519 597
rect 525 591 531 597
rect 537 591 543 597
rect 549 591 555 597
rect 561 591 567 597
rect 573 591 579 597
rect 585 591 591 597
rect 597 591 603 597
rect 609 591 615 597
rect 621 591 627 597
rect 633 591 639 597
rect 645 591 651 597
rect 657 591 663 597
rect 669 591 675 597
rect 681 591 687 597
rect 693 591 699 597
rect 705 591 711 597
rect 717 591 723 597
rect 729 591 735 597
rect 741 591 747 597
rect 753 591 759 597
rect 765 591 771 597
rect 777 591 783 597
rect 789 591 795 597
rect 801 591 807 597
rect 813 591 819 597
rect 825 591 831 597
rect 837 591 843 597
rect 849 591 855 597
rect 861 591 867 597
rect 873 591 879 597
rect 885 591 891 597
rect 897 591 903 597
rect 909 591 915 597
rect 921 591 927 597
rect 933 591 939 597
rect 945 591 951 597
rect 957 591 963 597
rect 969 591 975 597
rect 981 591 987 597
rect 993 591 999 597
rect 1005 591 1011 597
rect 1017 591 1023 597
rect 1029 591 1035 597
rect 1041 591 1047 597
rect 1053 591 1059 597
rect 1065 591 1071 597
rect 1077 591 1083 597
rect 1089 591 1095 597
rect 1101 591 1107 597
rect 1113 591 1119 597
rect 1125 591 1131 597
rect 1137 591 1143 597
rect 1149 591 1155 597
rect 1161 591 1167 597
rect 1173 591 1179 597
rect 1185 591 1191 597
rect 1197 591 1203 597
rect 1209 591 1215 597
rect 1221 591 1227 597
rect 1233 591 1239 597
rect 1245 591 1251 597
rect 1257 591 1263 597
rect 1269 591 1275 597
rect 1281 591 1287 597
rect 1293 591 1299 597
rect 1305 591 1311 597
rect 1317 591 1323 597
rect 1329 591 1335 597
rect 1341 591 1347 597
rect 1353 591 1359 597
rect 1365 591 1371 597
rect 1377 591 1383 597
rect 1389 591 1395 597
rect 1401 591 1407 597
rect 1413 591 1419 597
rect 1425 591 1431 597
rect 1437 591 1443 597
rect 1449 591 1455 597
rect 1461 591 1467 597
rect 1473 591 1479 597
rect 1485 591 1491 597
rect 1497 591 1503 597
rect 1509 591 1515 597
rect 1521 591 1527 597
rect 1533 591 1539 597
rect 1545 591 1551 597
rect 1557 591 1563 597
rect 1569 591 1575 597
rect 1581 591 1587 597
rect 1593 591 1599 597
rect 1605 591 1608 597
rect -84 588 1608 591
rect -84 585 -72 588
rect -84 579 -81 585
rect -75 579 -72 585
rect -84 573 -72 579
rect 1596 585 1608 588
rect 1596 579 1599 585
rect 1605 579 1608 585
rect -84 567 -81 573
rect -75 567 -72 573
rect -84 561 -72 567
rect -48 573 -12 576
rect -48 567 -45 573
rect -39 567 -33 573
rect -27 567 -21 573
rect -15 567 -12 573
rect -48 564 -12 567
rect 0 573 84 576
rect 0 567 3 573
rect 9 567 15 573
rect 21 567 27 573
rect 33 567 51 573
rect 57 567 63 573
rect 69 567 75 573
rect 81 567 84 573
rect 0 564 84 567
rect 96 573 180 576
rect 96 567 99 573
rect 105 567 111 573
rect 117 567 123 573
rect 129 567 147 573
rect 153 567 159 573
rect 165 567 171 573
rect 177 567 180 573
rect 96 564 180 567
rect 192 573 276 576
rect 192 567 195 573
rect 201 567 207 573
rect 213 567 219 573
rect 225 567 243 573
rect 249 567 255 573
rect 261 567 267 573
rect 273 567 276 573
rect 192 564 276 567
rect 288 573 372 576
rect 288 567 291 573
rect 297 567 303 573
rect 309 567 315 573
rect 321 567 339 573
rect 345 567 351 573
rect 357 567 363 573
rect 369 567 372 573
rect 288 564 372 567
rect 384 573 468 576
rect 384 567 387 573
rect 393 567 399 573
rect 405 567 411 573
rect 417 567 435 573
rect 441 567 447 573
rect 453 567 459 573
rect 465 567 468 573
rect 384 564 468 567
rect 480 573 564 576
rect 480 567 483 573
rect 489 567 495 573
rect 501 567 507 573
rect 513 567 531 573
rect 537 567 543 573
rect 549 567 555 573
rect 561 567 564 573
rect 480 564 564 567
rect 576 573 660 576
rect 576 567 579 573
rect 585 567 591 573
rect 597 567 603 573
rect 609 567 627 573
rect 633 567 639 573
rect 645 567 651 573
rect 657 567 660 573
rect 576 564 660 567
rect 672 573 756 576
rect 672 567 675 573
rect 681 567 687 573
rect 693 567 699 573
rect 705 567 723 573
rect 729 567 735 573
rect 741 567 747 573
rect 753 567 756 573
rect 672 564 756 567
rect 768 573 852 576
rect 768 567 771 573
rect 777 567 783 573
rect 789 567 795 573
rect 801 567 819 573
rect 825 567 831 573
rect 837 567 843 573
rect 849 567 852 573
rect 768 564 852 567
rect 864 573 948 576
rect 864 567 867 573
rect 873 567 879 573
rect 885 567 891 573
rect 897 567 915 573
rect 921 567 927 573
rect 933 567 939 573
rect 945 567 948 573
rect 864 564 948 567
rect 960 573 1044 576
rect 960 567 963 573
rect 969 567 975 573
rect 981 567 987 573
rect 993 567 1011 573
rect 1017 567 1023 573
rect 1029 567 1035 573
rect 1041 567 1044 573
rect 960 564 1044 567
rect 1056 573 1140 576
rect 1056 567 1059 573
rect 1065 567 1071 573
rect 1077 567 1083 573
rect 1089 567 1107 573
rect 1113 567 1119 573
rect 1125 567 1131 573
rect 1137 567 1140 573
rect 1056 564 1140 567
rect 1152 573 1236 576
rect 1152 567 1155 573
rect 1161 567 1167 573
rect 1173 567 1179 573
rect 1185 567 1203 573
rect 1209 567 1215 573
rect 1221 567 1227 573
rect 1233 567 1236 573
rect 1152 564 1236 567
rect 1248 573 1332 576
rect 1248 567 1251 573
rect 1257 567 1263 573
rect 1269 567 1275 573
rect 1281 567 1299 573
rect 1305 567 1311 573
rect 1317 567 1323 573
rect 1329 567 1332 573
rect 1248 564 1332 567
rect 1344 573 1428 576
rect 1344 567 1347 573
rect 1353 567 1359 573
rect 1365 567 1371 573
rect 1377 567 1395 573
rect 1401 567 1407 573
rect 1413 567 1419 573
rect 1425 567 1428 573
rect 1344 564 1428 567
rect 1440 573 1524 576
rect 1440 567 1443 573
rect 1449 567 1455 573
rect 1461 567 1467 573
rect 1473 567 1491 573
rect 1497 567 1503 573
rect 1509 567 1515 573
rect 1521 567 1524 573
rect 1440 564 1524 567
rect 1536 573 1572 576
rect 1536 567 1539 573
rect 1545 567 1551 573
rect 1557 567 1563 573
rect 1569 567 1572 573
rect 1536 564 1572 567
rect 1596 573 1608 579
rect 1596 567 1599 573
rect 1605 567 1608 573
rect -84 555 -81 561
rect -75 555 -72 561
rect -84 549 -72 555
rect 1596 561 1608 567
rect 1596 555 1599 561
rect 1605 555 1608 561
rect -84 543 -81 549
rect -75 543 -72 549
rect -84 537 -72 543
rect -84 531 -81 537
rect -75 531 -72 537
rect -84 525 -72 531
rect -84 519 -81 525
rect -75 519 -72 525
rect -84 513 -72 519
rect -60 549 -48 552
rect -60 543 -57 549
rect -51 543 -48 549
rect -60 537 -48 543
rect -60 531 -57 537
rect -51 531 -48 537
rect -60 525 -48 531
rect -60 519 -57 525
rect -51 519 -48 525
rect -60 516 -48 519
rect -36 549 -24 552
rect -36 543 -33 549
rect -27 543 -24 549
rect -36 537 -24 543
rect -36 531 -33 537
rect -27 531 -24 537
rect -36 525 -24 531
rect -36 519 -33 525
rect -27 519 -24 525
rect -84 507 -81 513
rect -75 507 -72 513
rect -84 504 -72 507
rect -36 504 -24 519
rect -12 549 0 552
rect -12 543 -9 549
rect -3 543 0 549
rect -12 537 0 543
rect -12 531 -9 537
rect -3 531 0 537
rect -12 525 0 531
rect -12 519 -9 525
rect -3 519 0 525
rect -12 516 0 519
rect 12 549 24 552
rect 12 543 15 549
rect 21 543 24 549
rect 12 537 24 543
rect 12 531 15 537
rect 21 531 24 537
rect 12 525 24 531
rect 12 519 15 525
rect 21 519 24 525
rect 12 504 24 519
rect 36 549 48 552
rect 36 543 39 549
rect 45 543 48 549
rect 36 537 48 543
rect 36 531 39 537
rect 45 531 48 537
rect 36 525 48 531
rect 36 519 39 525
rect 45 519 48 525
rect 36 516 48 519
rect 60 549 72 552
rect 60 543 63 549
rect 69 543 72 549
rect 60 537 72 543
rect 60 531 63 537
rect 69 531 72 537
rect 60 525 72 531
rect 60 519 63 525
rect 69 519 72 525
rect 60 504 72 519
rect 84 549 96 552
rect 84 543 87 549
rect 93 543 96 549
rect 84 537 96 543
rect 84 531 87 537
rect 93 531 96 537
rect 84 525 96 531
rect 84 519 87 525
rect 93 519 96 525
rect 84 516 96 519
rect 108 549 120 552
rect 108 543 111 549
rect 117 543 120 549
rect 108 537 120 543
rect 108 531 111 537
rect 117 531 120 537
rect 108 525 120 531
rect 108 519 111 525
rect 117 519 120 525
rect 108 504 120 519
rect 132 549 144 552
rect 132 543 135 549
rect 141 543 144 549
rect 132 537 144 543
rect 132 531 135 537
rect 141 531 144 537
rect 132 525 144 531
rect 132 519 135 525
rect 141 519 144 525
rect 132 516 144 519
rect 156 549 168 552
rect 156 543 159 549
rect 165 543 168 549
rect 156 537 168 543
rect 156 531 159 537
rect 165 531 168 537
rect 156 525 168 531
rect 156 519 159 525
rect 165 519 168 525
rect 156 504 168 519
rect 180 549 192 552
rect 180 543 183 549
rect 189 543 192 549
rect 180 537 192 543
rect 180 531 183 537
rect 189 531 192 537
rect 180 525 192 531
rect 180 519 183 525
rect 189 519 192 525
rect 180 516 192 519
rect 204 549 216 552
rect 204 543 207 549
rect 213 543 216 549
rect 204 537 216 543
rect 204 531 207 537
rect 213 531 216 537
rect 204 525 216 531
rect 204 519 207 525
rect 213 519 216 525
rect 204 504 216 519
rect 228 549 240 552
rect 228 543 231 549
rect 237 543 240 549
rect 228 537 240 543
rect 228 531 231 537
rect 237 531 240 537
rect 228 525 240 531
rect 228 519 231 525
rect 237 519 240 525
rect 228 516 240 519
rect 252 549 264 552
rect 252 543 255 549
rect 261 543 264 549
rect 252 537 264 543
rect 252 531 255 537
rect 261 531 264 537
rect 252 525 264 531
rect 252 519 255 525
rect 261 519 264 525
rect 252 504 264 519
rect 276 549 288 552
rect 276 543 279 549
rect 285 543 288 549
rect 276 537 288 543
rect 276 531 279 537
rect 285 531 288 537
rect 276 525 288 531
rect 276 519 279 525
rect 285 519 288 525
rect 276 516 288 519
rect 300 549 312 552
rect 300 543 303 549
rect 309 543 312 549
rect 300 537 312 543
rect 300 531 303 537
rect 309 531 312 537
rect 300 525 312 531
rect 300 519 303 525
rect 309 519 312 525
rect 300 504 312 519
rect 324 549 336 552
rect 324 543 327 549
rect 333 543 336 549
rect 324 537 336 543
rect 324 531 327 537
rect 333 531 336 537
rect 324 525 336 531
rect 324 519 327 525
rect 333 519 336 525
rect 324 516 336 519
rect 348 549 360 552
rect 348 543 351 549
rect 357 543 360 549
rect 348 537 360 543
rect 348 531 351 537
rect 357 531 360 537
rect 348 525 360 531
rect 348 519 351 525
rect 357 519 360 525
rect 348 504 360 519
rect 372 549 384 552
rect 372 543 375 549
rect 381 543 384 549
rect 372 537 384 543
rect 372 531 375 537
rect 381 531 384 537
rect 372 525 384 531
rect 372 519 375 525
rect 381 519 384 525
rect 372 516 384 519
rect 396 549 408 552
rect 396 543 399 549
rect 405 543 408 549
rect 396 537 408 543
rect 396 531 399 537
rect 405 531 408 537
rect 396 525 408 531
rect 396 519 399 525
rect 405 519 408 525
rect 396 504 408 519
rect 420 549 432 552
rect 420 543 423 549
rect 429 543 432 549
rect 420 537 432 543
rect 420 531 423 537
rect 429 531 432 537
rect 420 525 432 531
rect 420 519 423 525
rect 429 519 432 525
rect 420 516 432 519
rect 444 549 456 552
rect 444 543 447 549
rect 453 543 456 549
rect 444 537 456 543
rect 444 531 447 537
rect 453 531 456 537
rect 444 525 456 531
rect 444 519 447 525
rect 453 519 456 525
rect 444 504 456 519
rect 468 549 480 552
rect 468 543 471 549
rect 477 543 480 549
rect 468 537 480 543
rect 468 531 471 537
rect 477 531 480 537
rect 468 525 480 531
rect 468 519 471 525
rect 477 519 480 525
rect 468 516 480 519
rect 492 549 504 552
rect 492 543 495 549
rect 501 543 504 549
rect 492 537 504 543
rect 492 531 495 537
rect 501 531 504 537
rect 492 525 504 531
rect 492 519 495 525
rect 501 519 504 525
rect 492 504 504 519
rect 516 549 528 552
rect 516 543 519 549
rect 525 543 528 549
rect 516 537 528 543
rect 516 531 519 537
rect 525 531 528 537
rect 516 525 528 531
rect 516 519 519 525
rect 525 519 528 525
rect 516 516 528 519
rect 540 549 552 552
rect 540 543 543 549
rect 549 543 552 549
rect 540 537 552 543
rect 540 531 543 537
rect 549 531 552 537
rect 540 525 552 531
rect 540 519 543 525
rect 549 519 552 525
rect 540 504 552 519
rect 564 549 576 552
rect 564 543 567 549
rect 573 543 576 549
rect 564 537 576 543
rect 564 531 567 537
rect 573 531 576 537
rect 564 525 576 531
rect 564 519 567 525
rect 573 519 576 525
rect 564 516 576 519
rect 588 549 600 552
rect 588 543 591 549
rect 597 543 600 549
rect 588 537 600 543
rect 588 531 591 537
rect 597 531 600 537
rect 588 525 600 531
rect 588 519 591 525
rect 597 519 600 525
rect 588 504 600 519
rect 612 549 624 552
rect 612 543 615 549
rect 621 543 624 549
rect 612 537 624 543
rect 612 531 615 537
rect 621 531 624 537
rect 612 525 624 531
rect 612 519 615 525
rect 621 519 624 525
rect 612 516 624 519
rect 636 549 648 552
rect 636 543 639 549
rect 645 543 648 549
rect 636 537 648 543
rect 636 531 639 537
rect 645 531 648 537
rect 636 525 648 531
rect 636 519 639 525
rect 645 519 648 525
rect 636 504 648 519
rect 660 549 672 552
rect 660 543 663 549
rect 669 543 672 549
rect 660 537 672 543
rect 660 531 663 537
rect 669 531 672 537
rect 660 525 672 531
rect 660 519 663 525
rect 669 519 672 525
rect 660 516 672 519
rect 684 549 696 552
rect 684 543 687 549
rect 693 543 696 549
rect 684 537 696 543
rect 684 531 687 537
rect 693 531 696 537
rect 684 525 696 531
rect 684 519 687 525
rect 693 519 696 525
rect 684 504 696 519
rect 708 549 720 552
rect 708 543 711 549
rect 717 543 720 549
rect 708 537 720 543
rect 708 531 711 537
rect 717 531 720 537
rect 708 525 720 531
rect 708 519 711 525
rect 717 519 720 525
rect 708 516 720 519
rect 732 549 744 552
rect 732 543 735 549
rect 741 543 744 549
rect 732 537 744 543
rect 732 531 735 537
rect 741 531 744 537
rect 732 525 744 531
rect 732 519 735 525
rect 741 519 744 525
rect 732 504 744 519
rect 756 549 768 552
rect 756 543 759 549
rect 765 543 768 549
rect 756 537 768 543
rect 756 531 759 537
rect 765 531 768 537
rect 756 525 768 531
rect 756 519 759 525
rect 765 519 768 525
rect 756 516 768 519
rect 780 549 792 552
rect 780 543 783 549
rect 789 543 792 549
rect 780 537 792 543
rect 780 531 783 537
rect 789 531 792 537
rect 780 525 792 531
rect 780 519 783 525
rect 789 519 792 525
rect 780 504 792 519
rect 804 549 816 552
rect 804 543 807 549
rect 813 543 816 549
rect 804 537 816 543
rect 804 531 807 537
rect 813 531 816 537
rect 804 525 816 531
rect 804 519 807 525
rect 813 519 816 525
rect 804 516 816 519
rect 828 549 840 552
rect 828 543 831 549
rect 837 543 840 549
rect 828 537 840 543
rect 828 531 831 537
rect 837 531 840 537
rect 828 525 840 531
rect 828 519 831 525
rect 837 519 840 525
rect 828 504 840 519
rect 852 549 864 552
rect 852 543 855 549
rect 861 543 864 549
rect 852 537 864 543
rect 852 531 855 537
rect 861 531 864 537
rect 852 525 864 531
rect 852 519 855 525
rect 861 519 864 525
rect 852 516 864 519
rect 876 549 888 552
rect 876 543 879 549
rect 885 543 888 549
rect 876 537 888 543
rect 876 531 879 537
rect 885 531 888 537
rect 876 525 888 531
rect 876 519 879 525
rect 885 519 888 525
rect 876 504 888 519
rect 900 549 912 552
rect 900 543 903 549
rect 909 543 912 549
rect 900 537 912 543
rect 900 531 903 537
rect 909 531 912 537
rect 900 525 912 531
rect 900 519 903 525
rect 909 519 912 525
rect 900 516 912 519
rect 924 549 936 552
rect 924 543 927 549
rect 933 543 936 549
rect 924 537 936 543
rect 924 531 927 537
rect 933 531 936 537
rect 924 525 936 531
rect 924 519 927 525
rect 933 519 936 525
rect 924 504 936 519
rect 948 549 960 552
rect 948 543 951 549
rect 957 543 960 549
rect 948 537 960 543
rect 948 531 951 537
rect 957 531 960 537
rect 948 525 960 531
rect 948 519 951 525
rect 957 519 960 525
rect 948 516 960 519
rect 972 549 984 552
rect 972 543 975 549
rect 981 543 984 549
rect 972 537 984 543
rect 972 531 975 537
rect 981 531 984 537
rect 972 525 984 531
rect 972 519 975 525
rect 981 519 984 525
rect 972 504 984 519
rect 996 549 1008 552
rect 996 543 999 549
rect 1005 543 1008 549
rect 996 537 1008 543
rect 996 531 999 537
rect 1005 531 1008 537
rect 996 525 1008 531
rect 996 519 999 525
rect 1005 519 1008 525
rect 996 516 1008 519
rect 1020 549 1032 552
rect 1020 543 1023 549
rect 1029 543 1032 549
rect 1020 537 1032 543
rect 1020 531 1023 537
rect 1029 531 1032 537
rect 1020 525 1032 531
rect 1020 519 1023 525
rect 1029 519 1032 525
rect 1020 504 1032 519
rect 1044 549 1056 552
rect 1044 543 1047 549
rect 1053 543 1056 549
rect 1044 537 1056 543
rect 1044 531 1047 537
rect 1053 531 1056 537
rect 1044 525 1056 531
rect 1044 519 1047 525
rect 1053 519 1056 525
rect 1044 516 1056 519
rect 1068 549 1080 552
rect 1068 543 1071 549
rect 1077 543 1080 549
rect 1068 537 1080 543
rect 1068 531 1071 537
rect 1077 531 1080 537
rect 1068 525 1080 531
rect 1068 519 1071 525
rect 1077 519 1080 525
rect 1068 504 1080 519
rect 1092 549 1104 552
rect 1092 543 1095 549
rect 1101 543 1104 549
rect 1092 537 1104 543
rect 1092 531 1095 537
rect 1101 531 1104 537
rect 1092 525 1104 531
rect 1092 519 1095 525
rect 1101 519 1104 525
rect 1092 516 1104 519
rect 1116 549 1128 552
rect 1116 543 1119 549
rect 1125 543 1128 549
rect 1116 537 1128 543
rect 1116 531 1119 537
rect 1125 531 1128 537
rect 1116 525 1128 531
rect 1116 519 1119 525
rect 1125 519 1128 525
rect 1116 504 1128 519
rect 1140 549 1152 552
rect 1140 543 1143 549
rect 1149 543 1152 549
rect 1140 537 1152 543
rect 1140 531 1143 537
rect 1149 531 1152 537
rect 1140 525 1152 531
rect 1140 519 1143 525
rect 1149 519 1152 525
rect 1140 516 1152 519
rect 1164 549 1176 552
rect 1164 543 1167 549
rect 1173 543 1176 549
rect 1164 537 1176 543
rect 1164 531 1167 537
rect 1173 531 1176 537
rect 1164 525 1176 531
rect 1164 519 1167 525
rect 1173 519 1176 525
rect 1164 504 1176 519
rect 1188 549 1200 552
rect 1188 543 1191 549
rect 1197 543 1200 549
rect 1188 537 1200 543
rect 1188 531 1191 537
rect 1197 531 1200 537
rect 1188 525 1200 531
rect 1188 519 1191 525
rect 1197 519 1200 525
rect 1188 516 1200 519
rect 1212 549 1224 552
rect 1212 543 1215 549
rect 1221 543 1224 549
rect 1212 537 1224 543
rect 1212 531 1215 537
rect 1221 531 1224 537
rect 1212 525 1224 531
rect 1212 519 1215 525
rect 1221 519 1224 525
rect 1212 504 1224 519
rect 1236 549 1248 552
rect 1236 543 1239 549
rect 1245 543 1248 549
rect 1236 537 1248 543
rect 1236 531 1239 537
rect 1245 531 1248 537
rect 1236 525 1248 531
rect 1236 519 1239 525
rect 1245 519 1248 525
rect 1236 516 1248 519
rect 1260 549 1272 552
rect 1260 543 1263 549
rect 1269 543 1272 549
rect 1260 537 1272 543
rect 1260 531 1263 537
rect 1269 531 1272 537
rect 1260 525 1272 531
rect 1260 519 1263 525
rect 1269 519 1272 525
rect 1260 504 1272 519
rect 1284 549 1296 552
rect 1284 543 1287 549
rect 1293 543 1296 549
rect 1284 537 1296 543
rect 1284 531 1287 537
rect 1293 531 1296 537
rect 1284 525 1296 531
rect 1284 519 1287 525
rect 1293 519 1296 525
rect 1284 516 1296 519
rect 1308 549 1320 552
rect 1308 543 1311 549
rect 1317 543 1320 549
rect 1308 537 1320 543
rect 1308 531 1311 537
rect 1317 531 1320 537
rect 1308 525 1320 531
rect 1308 519 1311 525
rect 1317 519 1320 525
rect 1308 504 1320 519
rect 1332 549 1344 552
rect 1332 543 1335 549
rect 1341 543 1344 549
rect 1332 537 1344 543
rect 1332 531 1335 537
rect 1341 531 1344 537
rect 1332 525 1344 531
rect 1332 519 1335 525
rect 1341 519 1344 525
rect 1332 516 1344 519
rect 1356 549 1368 552
rect 1356 543 1359 549
rect 1365 543 1368 549
rect 1356 537 1368 543
rect 1356 531 1359 537
rect 1365 531 1368 537
rect 1356 525 1368 531
rect 1356 519 1359 525
rect 1365 519 1368 525
rect 1356 504 1368 519
rect 1380 549 1392 552
rect 1380 543 1383 549
rect 1389 543 1392 549
rect 1380 537 1392 543
rect 1380 531 1383 537
rect 1389 531 1392 537
rect 1380 525 1392 531
rect 1380 519 1383 525
rect 1389 519 1392 525
rect 1380 516 1392 519
rect 1404 549 1416 552
rect 1404 543 1407 549
rect 1413 543 1416 549
rect 1404 537 1416 543
rect 1404 531 1407 537
rect 1413 531 1416 537
rect 1404 525 1416 531
rect 1404 519 1407 525
rect 1413 519 1416 525
rect 1404 504 1416 519
rect 1428 549 1440 552
rect 1428 543 1431 549
rect 1437 543 1440 549
rect 1428 537 1440 543
rect 1428 531 1431 537
rect 1437 531 1440 537
rect 1428 525 1440 531
rect 1428 519 1431 525
rect 1437 519 1440 525
rect 1428 516 1440 519
rect 1452 549 1464 552
rect 1452 543 1455 549
rect 1461 543 1464 549
rect 1452 537 1464 543
rect 1452 531 1455 537
rect 1461 531 1464 537
rect 1452 525 1464 531
rect 1452 519 1455 525
rect 1461 519 1464 525
rect 1452 504 1464 519
rect 1476 549 1488 552
rect 1476 543 1479 549
rect 1485 543 1488 549
rect 1476 537 1488 543
rect 1476 531 1479 537
rect 1485 531 1488 537
rect 1476 525 1488 531
rect 1476 519 1479 525
rect 1485 519 1488 525
rect 1476 516 1488 519
rect 1500 549 1512 552
rect 1500 543 1503 549
rect 1509 543 1512 549
rect 1500 537 1512 543
rect 1500 531 1503 537
rect 1509 531 1512 537
rect 1500 525 1512 531
rect 1500 519 1503 525
rect 1509 519 1512 525
rect 1500 504 1512 519
rect 1524 549 1536 552
rect 1524 543 1527 549
rect 1533 543 1536 549
rect 1524 537 1536 543
rect 1524 531 1527 537
rect 1533 531 1536 537
rect 1524 525 1536 531
rect 1524 519 1527 525
rect 1533 519 1536 525
rect 1524 516 1536 519
rect 1548 549 1560 552
rect 1548 543 1551 549
rect 1557 543 1560 549
rect 1548 537 1560 543
rect 1548 531 1551 537
rect 1557 531 1560 537
rect 1548 525 1560 531
rect 1548 519 1551 525
rect 1557 519 1560 525
rect 1548 504 1560 519
rect 1572 549 1584 552
rect 1572 543 1575 549
rect 1581 543 1584 549
rect 1572 537 1584 543
rect 1572 531 1575 537
rect 1581 531 1584 537
rect 1572 525 1584 531
rect 1572 519 1575 525
rect 1581 519 1584 525
rect 1572 516 1584 519
rect 1596 549 1608 555
rect 1596 543 1599 549
rect 1605 543 1608 549
rect 1596 537 1608 543
rect 1596 531 1599 537
rect 1605 531 1608 537
rect 1596 525 1608 531
rect 1596 519 1599 525
rect 1605 519 1608 525
rect 1596 513 1608 519
rect 1596 507 1599 513
rect 1605 507 1608 513
rect 1596 504 1608 507
rect -84 501 1608 504
rect -84 495 -81 501
rect -75 495 -69 501
rect -63 495 -57 501
rect -51 495 -45 501
rect -39 495 -33 501
rect -27 495 -21 501
rect -15 495 -9 501
rect -3 495 3 501
rect 9 495 15 501
rect 21 495 27 501
rect 33 495 39 501
rect 45 495 51 501
rect 57 495 63 501
rect 69 495 75 501
rect 81 495 87 501
rect 93 495 99 501
rect 105 495 111 501
rect 117 495 123 501
rect 129 495 135 501
rect 141 495 147 501
rect 153 495 159 501
rect 165 495 171 501
rect 177 495 183 501
rect 189 495 195 501
rect 201 495 207 501
rect 213 495 219 501
rect 225 495 231 501
rect 237 495 243 501
rect 249 495 255 501
rect 261 495 267 501
rect 273 495 279 501
rect 285 495 291 501
rect 297 495 303 501
rect 309 495 315 501
rect 321 495 327 501
rect 333 495 339 501
rect 345 495 351 501
rect 357 495 363 501
rect 369 495 375 501
rect 381 495 387 501
rect 393 495 399 501
rect 405 495 411 501
rect 417 495 423 501
rect 429 495 435 501
rect 441 495 447 501
rect 453 495 459 501
rect 465 495 471 501
rect 477 495 483 501
rect 489 495 495 501
rect 501 495 507 501
rect 513 495 519 501
rect 525 495 531 501
rect 537 495 543 501
rect 549 495 555 501
rect 561 495 567 501
rect 573 495 579 501
rect 585 495 591 501
rect 597 495 603 501
rect 609 495 615 501
rect 621 495 627 501
rect 633 495 639 501
rect 645 495 651 501
rect 657 495 663 501
rect 669 495 675 501
rect 681 495 687 501
rect 693 495 699 501
rect 705 495 711 501
rect 717 495 723 501
rect 729 495 735 501
rect 741 495 747 501
rect 753 495 759 501
rect 765 495 771 501
rect 777 495 783 501
rect 789 495 795 501
rect 801 495 807 501
rect 813 495 819 501
rect 825 495 831 501
rect 837 495 843 501
rect 849 495 855 501
rect 861 495 867 501
rect 873 495 879 501
rect 885 495 891 501
rect 897 495 903 501
rect 909 495 915 501
rect 921 495 927 501
rect 933 495 939 501
rect 945 495 951 501
rect 957 495 963 501
rect 969 495 975 501
rect 981 495 987 501
rect 993 495 999 501
rect 1005 495 1011 501
rect 1017 495 1023 501
rect 1029 495 1035 501
rect 1041 495 1047 501
rect 1053 495 1059 501
rect 1065 495 1071 501
rect 1077 495 1083 501
rect 1089 495 1095 501
rect 1101 495 1107 501
rect 1113 495 1119 501
rect 1125 495 1131 501
rect 1137 495 1143 501
rect 1149 495 1155 501
rect 1161 495 1167 501
rect 1173 495 1179 501
rect 1185 495 1191 501
rect 1197 495 1203 501
rect 1209 495 1215 501
rect 1221 495 1227 501
rect 1233 495 1239 501
rect 1245 495 1251 501
rect 1257 495 1263 501
rect 1269 495 1275 501
rect 1281 495 1287 501
rect 1293 495 1299 501
rect 1305 495 1311 501
rect 1317 495 1323 501
rect 1329 495 1335 501
rect 1341 495 1347 501
rect 1353 495 1359 501
rect 1365 495 1371 501
rect 1377 495 1383 501
rect 1389 495 1395 501
rect 1401 495 1407 501
rect 1413 495 1419 501
rect 1425 495 1431 501
rect 1437 495 1443 501
rect 1449 495 1455 501
rect 1461 495 1467 501
rect 1473 495 1479 501
rect 1485 495 1491 501
rect 1497 495 1503 501
rect 1509 495 1515 501
rect 1521 495 1527 501
rect 1533 495 1539 501
rect 1545 495 1551 501
rect 1557 495 1563 501
rect 1569 495 1575 501
rect 1581 495 1587 501
rect 1593 495 1599 501
rect 1605 495 1608 501
rect -84 492 1608 495
rect 1620 597 1632 603
rect 1620 591 1623 597
rect 1629 591 1632 597
rect 1620 585 1632 591
rect 1620 579 1623 585
rect 1629 579 1632 585
rect 1620 573 1632 579
rect 1620 567 1623 573
rect 1629 567 1632 573
rect 1620 561 1632 567
rect 1620 555 1623 561
rect 1629 555 1632 561
rect 1620 549 1632 555
rect 1620 543 1623 549
rect 1629 543 1632 549
rect 1620 537 1632 543
rect 1620 531 1623 537
rect 1629 531 1632 537
rect 1620 525 1632 531
rect 1620 519 1623 525
rect 1629 519 1632 525
rect 1620 513 1632 519
rect 1620 507 1623 513
rect 1629 507 1632 513
rect 1620 501 1632 507
rect 1620 495 1623 501
rect 1629 495 1632 501
rect -108 483 -105 489
rect -99 483 -96 489
rect -108 480 -96 483
rect 1620 489 1632 495
rect 1620 483 1623 489
rect 1629 483 1632 489
rect 1620 480 1632 483
rect -108 477 1632 480
rect -108 471 -105 477
rect -99 471 -93 477
rect -87 471 -81 477
rect -75 471 -69 477
rect -63 471 -57 477
rect -51 471 -45 477
rect -39 471 -33 477
rect -27 471 -21 477
rect -15 471 -9 477
rect -3 471 3 477
rect 9 471 15 477
rect 21 471 27 477
rect 33 471 39 477
rect 45 471 51 477
rect 57 471 63 477
rect 69 471 75 477
rect 81 471 87 477
rect 93 471 99 477
rect 105 471 111 477
rect 117 471 123 477
rect 129 471 135 477
rect 141 471 147 477
rect 153 471 159 477
rect 165 471 171 477
rect 177 471 183 477
rect 189 471 195 477
rect 201 471 207 477
rect 213 471 219 477
rect 225 471 231 477
rect 237 471 243 477
rect 249 471 255 477
rect 261 471 267 477
rect 273 471 279 477
rect 285 471 291 477
rect 297 471 303 477
rect 309 471 315 477
rect 321 471 327 477
rect 333 471 339 477
rect 345 471 351 477
rect 357 471 363 477
rect 369 471 375 477
rect 381 471 387 477
rect 393 471 399 477
rect 405 471 411 477
rect 417 471 423 477
rect 429 471 435 477
rect 441 471 447 477
rect 453 471 459 477
rect 465 471 471 477
rect 477 471 483 477
rect 489 471 495 477
rect 501 471 507 477
rect 513 471 519 477
rect 525 471 531 477
rect 537 471 543 477
rect 549 471 555 477
rect 561 471 567 477
rect 573 471 579 477
rect 585 471 591 477
rect 597 471 603 477
rect 609 471 615 477
rect 621 471 627 477
rect 633 471 639 477
rect 645 471 651 477
rect 657 471 663 477
rect 669 471 675 477
rect 681 471 687 477
rect 693 471 699 477
rect 705 471 711 477
rect 717 471 723 477
rect 729 471 735 477
rect 741 471 747 477
rect 753 471 759 477
rect 765 471 771 477
rect 777 471 783 477
rect 789 471 795 477
rect 801 471 807 477
rect 813 471 819 477
rect 825 471 831 477
rect 837 471 843 477
rect 849 471 855 477
rect 861 471 867 477
rect 873 471 879 477
rect 885 471 891 477
rect 897 471 903 477
rect 909 471 915 477
rect 921 471 927 477
rect 933 471 939 477
rect 945 471 951 477
rect 957 471 963 477
rect 969 471 975 477
rect 981 471 987 477
rect 993 471 999 477
rect 1005 471 1011 477
rect 1017 471 1023 477
rect 1029 471 1035 477
rect 1041 471 1047 477
rect 1053 471 1059 477
rect 1065 471 1071 477
rect 1077 471 1083 477
rect 1089 471 1095 477
rect 1101 471 1107 477
rect 1113 471 1119 477
rect 1125 471 1131 477
rect 1137 471 1143 477
rect 1149 471 1155 477
rect 1161 471 1167 477
rect 1173 471 1179 477
rect 1185 471 1191 477
rect 1197 471 1203 477
rect 1209 471 1215 477
rect 1221 471 1227 477
rect 1233 471 1239 477
rect 1245 471 1251 477
rect 1257 471 1263 477
rect 1269 471 1275 477
rect 1281 471 1287 477
rect 1293 471 1299 477
rect 1305 471 1311 477
rect 1317 471 1323 477
rect 1329 471 1335 477
rect 1341 471 1347 477
rect 1353 471 1359 477
rect 1365 471 1371 477
rect 1377 471 1383 477
rect 1389 471 1395 477
rect 1401 471 1407 477
rect 1413 471 1419 477
rect 1425 471 1431 477
rect 1437 471 1443 477
rect 1449 471 1455 477
rect 1461 471 1467 477
rect 1473 471 1479 477
rect 1485 471 1491 477
rect 1497 471 1503 477
rect 1509 471 1515 477
rect 1521 471 1527 477
rect 1533 471 1539 477
rect 1545 471 1551 477
rect 1557 471 1563 477
rect 1569 471 1575 477
rect 1581 471 1587 477
rect 1593 471 1599 477
rect 1605 471 1611 477
rect 1617 471 1623 477
rect 1629 471 1632 477
rect -108 468 1632 471
rect -108 465 -96 468
rect -108 459 -105 465
rect -99 459 -96 465
rect -108 453 -96 459
rect 1620 465 1632 468
rect 1620 459 1623 465
rect 1629 459 1632 465
rect -108 447 -105 453
rect -99 447 -96 453
rect -108 441 -96 447
rect -108 435 -105 441
rect -99 435 -96 441
rect -108 429 -96 435
rect -108 423 -105 429
rect -99 423 -96 429
rect -108 417 -96 423
rect -108 411 -105 417
rect -99 411 -96 417
rect -108 405 -96 411
rect -108 399 -105 405
rect -99 399 -96 405
rect -108 393 -96 399
rect -108 387 -105 393
rect -99 387 -96 393
rect -108 381 -96 387
rect -108 375 -105 381
rect -99 375 -96 381
rect -108 369 -96 375
rect -108 363 -105 369
rect -99 363 -96 369
rect -108 357 -96 363
rect -108 351 -105 357
rect -99 351 -96 357
rect -108 345 -96 351
rect -84 453 1608 456
rect -84 447 -81 453
rect -75 447 -69 453
rect -63 447 -57 453
rect -51 447 -45 453
rect -39 447 -33 453
rect -27 447 -21 453
rect -15 447 -9 453
rect -3 447 3 453
rect 9 447 15 453
rect 21 447 27 453
rect 33 447 39 453
rect 45 447 51 453
rect 57 447 63 453
rect 69 447 75 453
rect 81 447 87 453
rect 93 447 99 453
rect 105 447 111 453
rect 117 447 123 453
rect 129 447 135 453
rect 141 447 147 453
rect 153 447 159 453
rect 165 447 171 453
rect 177 447 183 453
rect 189 447 195 453
rect 201 447 207 453
rect 213 447 219 453
rect 225 447 231 453
rect 237 447 243 453
rect 249 447 255 453
rect 261 447 267 453
rect 273 447 279 453
rect 285 447 291 453
rect 297 447 303 453
rect 309 447 315 453
rect 321 447 327 453
rect 333 447 339 453
rect 345 447 351 453
rect 357 447 363 453
rect 369 447 375 453
rect 381 447 387 453
rect 393 447 399 453
rect 405 447 411 453
rect 417 447 423 453
rect 429 447 435 453
rect 441 447 447 453
rect 453 447 459 453
rect 465 447 471 453
rect 477 447 483 453
rect 489 447 495 453
rect 501 447 507 453
rect 513 447 519 453
rect 525 447 531 453
rect 537 447 543 453
rect 549 447 555 453
rect 561 447 567 453
rect 573 447 579 453
rect 585 447 591 453
rect 597 447 603 453
rect 609 447 615 453
rect 621 447 627 453
rect 633 447 639 453
rect 645 447 651 453
rect 657 447 663 453
rect 669 447 675 453
rect 681 447 687 453
rect 693 447 699 453
rect 705 447 711 453
rect 717 447 723 453
rect 729 447 735 453
rect 741 447 747 453
rect 753 447 759 453
rect 765 447 771 453
rect 777 447 783 453
rect 789 447 795 453
rect 801 447 807 453
rect 813 447 819 453
rect 825 447 831 453
rect 837 447 843 453
rect 849 447 855 453
rect 861 447 867 453
rect 873 447 879 453
rect 885 447 891 453
rect 897 447 903 453
rect 909 447 915 453
rect 921 447 927 453
rect 933 447 939 453
rect 945 447 951 453
rect 957 447 963 453
rect 969 447 975 453
rect 981 447 987 453
rect 993 447 999 453
rect 1005 447 1011 453
rect 1017 447 1023 453
rect 1029 447 1035 453
rect 1041 447 1047 453
rect 1053 447 1059 453
rect 1065 447 1071 453
rect 1077 447 1083 453
rect 1089 447 1095 453
rect 1101 447 1107 453
rect 1113 447 1119 453
rect 1125 447 1131 453
rect 1137 447 1143 453
rect 1149 447 1155 453
rect 1161 447 1167 453
rect 1173 447 1179 453
rect 1185 447 1191 453
rect 1197 447 1203 453
rect 1209 447 1215 453
rect 1221 447 1227 453
rect 1233 447 1239 453
rect 1245 447 1251 453
rect 1257 447 1263 453
rect 1269 447 1275 453
rect 1281 447 1287 453
rect 1293 447 1299 453
rect 1305 447 1311 453
rect 1317 447 1323 453
rect 1329 447 1335 453
rect 1341 447 1347 453
rect 1353 447 1359 453
rect 1365 447 1371 453
rect 1377 447 1383 453
rect 1389 447 1395 453
rect 1401 447 1407 453
rect 1413 447 1419 453
rect 1425 447 1431 453
rect 1437 447 1443 453
rect 1449 447 1455 453
rect 1461 447 1467 453
rect 1473 447 1479 453
rect 1485 447 1491 453
rect 1497 447 1503 453
rect 1509 447 1515 453
rect 1521 447 1527 453
rect 1533 447 1539 453
rect 1545 447 1551 453
rect 1557 447 1563 453
rect 1569 447 1575 453
rect 1581 447 1587 453
rect 1593 447 1599 453
rect 1605 447 1608 453
rect -84 444 1608 447
rect -84 441 -72 444
rect -84 435 -81 441
rect -75 435 -72 441
rect -84 429 -72 435
rect 1596 441 1608 444
rect 1596 435 1599 441
rect 1605 435 1608 441
rect -84 423 -81 429
rect -75 423 -72 429
rect -84 417 -72 423
rect -84 411 -81 417
rect -75 411 -72 417
rect -84 405 -72 411
rect -84 399 -81 405
rect -75 399 -72 405
rect -84 393 -72 399
rect -60 429 -48 432
rect -60 423 -57 429
rect -51 423 -48 429
rect -60 417 -48 423
rect -12 429 0 432
rect -12 423 -9 429
rect -3 423 0 429
rect -60 411 -57 417
rect -51 411 -48 417
rect -60 405 -48 411
rect -60 399 -57 405
rect -51 399 -48 405
rect -60 396 -48 399
rect -36 417 -24 420
rect -36 411 -33 417
rect -27 411 -24 417
rect -36 405 -24 411
rect -36 399 -33 405
rect -27 399 -24 405
rect -84 387 -81 393
rect -75 387 -72 393
rect -84 381 -72 387
rect -36 384 -24 399
rect -12 417 0 423
rect 36 429 48 432
rect 36 423 39 429
rect 45 423 48 429
rect -12 411 -9 417
rect -3 411 0 417
rect -12 405 0 411
rect -12 399 -9 405
rect -3 399 0 405
rect -12 396 0 399
rect 12 417 24 420
rect 12 411 15 417
rect 21 411 24 417
rect 12 405 24 411
rect 12 399 15 405
rect 21 399 24 405
rect 12 396 24 399
rect 36 417 48 423
rect 84 429 96 432
rect 84 423 87 429
rect 93 423 96 429
rect 36 411 39 417
rect 45 411 48 417
rect 36 405 48 411
rect 36 399 39 405
rect 45 399 48 405
rect 36 396 48 399
rect 60 417 72 420
rect 60 411 63 417
rect 69 411 72 417
rect 60 405 72 411
rect 60 399 63 405
rect 69 399 72 405
rect 60 396 72 399
rect 84 417 96 423
rect 132 429 144 432
rect 132 423 135 429
rect 141 423 144 429
rect 84 411 87 417
rect 93 411 96 417
rect 84 405 96 411
rect 84 399 87 405
rect 93 399 96 405
rect 84 396 96 399
rect 108 417 120 420
rect 108 411 111 417
rect 117 411 120 417
rect 108 405 120 411
rect 108 399 111 405
rect 117 399 120 405
rect 108 396 120 399
rect 132 417 144 423
rect 180 429 192 432
rect 180 423 183 429
rect 189 423 192 429
rect 132 411 135 417
rect 141 411 144 417
rect 132 405 144 411
rect 132 399 135 405
rect 141 399 144 405
rect 132 396 144 399
rect 156 417 168 420
rect 156 411 159 417
rect 165 411 168 417
rect 156 405 168 411
rect 156 399 159 405
rect 165 399 168 405
rect 156 396 168 399
rect 180 417 192 423
rect 180 411 183 417
rect 189 411 192 417
rect 180 405 192 411
rect 180 399 183 405
rect 189 399 192 405
rect 180 396 192 399
rect 228 417 240 432
rect 228 411 231 417
rect 237 411 240 417
rect 228 405 240 411
rect 228 399 231 405
rect 237 399 240 405
rect 228 396 240 399
rect 276 429 288 432
rect 276 423 279 429
rect 285 423 288 429
rect 276 417 288 423
rect 276 411 279 417
rect 285 411 288 417
rect 276 405 288 411
rect 276 399 279 405
rect 285 399 288 405
rect 276 396 288 399
rect 324 417 336 432
rect 324 411 327 417
rect 333 411 336 417
rect 324 405 336 411
rect 324 399 327 405
rect 333 399 336 405
rect 324 396 336 399
rect 372 429 384 432
rect 372 423 375 429
rect 381 423 384 429
rect 372 417 384 423
rect 372 411 375 417
rect 381 411 384 417
rect 372 405 384 411
rect 372 399 375 405
rect 381 399 384 405
rect 372 396 384 399
rect 420 417 432 432
rect 420 411 423 417
rect 429 411 432 417
rect 420 405 432 411
rect 420 399 423 405
rect 429 399 432 405
rect 420 396 432 399
rect 468 429 480 432
rect 468 423 471 429
rect 477 423 480 429
rect 468 417 480 423
rect 468 411 471 417
rect 477 411 480 417
rect 468 405 480 411
rect 468 399 471 405
rect 477 399 480 405
rect 468 396 480 399
rect 516 417 528 432
rect 516 411 519 417
rect 525 411 528 417
rect 516 405 528 411
rect 516 399 519 405
rect 525 399 528 405
rect 516 396 528 399
rect 564 429 576 432
rect 564 423 567 429
rect 573 423 576 429
rect 564 417 576 423
rect 612 429 624 432
rect 612 423 615 429
rect 621 423 624 429
rect 564 411 567 417
rect 573 411 576 417
rect 564 405 576 411
rect 564 399 567 405
rect 573 399 576 405
rect 564 396 576 399
rect 588 417 600 420
rect 588 411 591 417
rect 597 411 600 417
rect 588 405 600 411
rect 588 399 591 405
rect 597 399 600 405
rect 588 396 600 399
rect 612 417 624 423
rect 660 429 672 432
rect 660 423 663 429
rect 669 423 672 429
rect 612 411 615 417
rect 621 411 624 417
rect 612 405 624 411
rect 612 399 615 405
rect 621 399 624 405
rect 612 396 624 399
rect 636 417 648 420
rect 636 411 639 417
rect 645 411 648 417
rect 636 405 648 411
rect 636 399 639 405
rect 645 399 648 405
rect 636 396 648 399
rect 660 417 672 423
rect 708 429 720 432
rect 708 423 711 429
rect 717 423 720 429
rect 660 411 663 417
rect 669 411 672 417
rect 660 405 672 411
rect 660 399 663 405
rect 669 399 672 405
rect 660 396 672 399
rect 684 417 696 420
rect 684 411 687 417
rect 693 411 696 417
rect 684 405 696 411
rect 684 399 687 405
rect 693 399 696 405
rect 684 396 696 399
rect 708 417 720 423
rect 756 429 768 432
rect 756 423 759 429
rect 765 423 768 429
rect 708 411 711 417
rect 717 411 720 417
rect 708 405 720 411
rect 708 399 711 405
rect 717 399 720 405
rect 708 396 720 399
rect 732 417 744 420
rect 732 411 735 417
rect 741 411 744 417
rect 732 405 744 411
rect 732 399 735 405
rect 741 399 744 405
rect 732 396 744 399
rect 756 417 768 423
rect 804 429 816 432
rect 804 423 807 429
rect 813 423 816 429
rect 756 411 759 417
rect 765 411 768 417
rect 756 405 768 411
rect 756 399 759 405
rect 765 399 768 405
rect 756 396 768 399
rect 780 417 792 420
rect 780 411 783 417
rect 789 411 792 417
rect 780 405 792 411
rect 780 399 783 405
rect 789 399 792 405
rect 780 396 792 399
rect 804 417 816 423
rect 852 429 864 432
rect 852 423 855 429
rect 861 423 864 429
rect 804 411 807 417
rect 813 411 816 417
rect 804 405 816 411
rect 804 399 807 405
rect 813 399 816 405
rect 804 396 816 399
rect 828 417 840 420
rect 828 411 831 417
rect 837 411 840 417
rect 828 405 840 411
rect 828 399 831 405
rect 837 399 840 405
rect 828 396 840 399
rect 852 417 864 423
rect 900 429 912 432
rect 900 423 903 429
rect 909 423 912 429
rect 852 411 855 417
rect 861 411 864 417
rect 852 405 864 411
rect 852 399 855 405
rect 861 399 864 405
rect 852 396 864 399
rect 876 417 888 420
rect 876 411 879 417
rect 885 411 888 417
rect 876 405 888 411
rect 876 399 879 405
rect 885 399 888 405
rect 876 396 888 399
rect 900 417 912 423
rect 948 429 960 432
rect 948 423 951 429
rect 957 423 960 429
rect 900 411 903 417
rect 909 411 912 417
rect 900 405 912 411
rect 900 399 903 405
rect 909 399 912 405
rect 900 396 912 399
rect 924 417 936 420
rect 924 411 927 417
rect 933 411 936 417
rect 924 405 936 411
rect 924 399 927 405
rect 933 399 936 405
rect 924 396 936 399
rect 948 417 960 423
rect 948 411 951 417
rect 957 411 960 417
rect 948 405 960 411
rect 948 399 951 405
rect 957 399 960 405
rect 948 396 960 399
rect 996 417 1008 432
rect 996 411 999 417
rect 1005 411 1008 417
rect 996 405 1008 411
rect 996 399 999 405
rect 1005 399 1008 405
rect 996 396 1008 399
rect 1044 429 1056 432
rect 1044 423 1047 429
rect 1053 423 1056 429
rect 1044 417 1056 423
rect 1044 411 1047 417
rect 1053 411 1056 417
rect 1044 405 1056 411
rect 1044 399 1047 405
rect 1053 399 1056 405
rect 1044 396 1056 399
rect 1092 417 1104 432
rect 1092 411 1095 417
rect 1101 411 1104 417
rect 1092 405 1104 411
rect 1092 399 1095 405
rect 1101 399 1104 405
rect 1092 396 1104 399
rect 1140 429 1152 432
rect 1140 423 1143 429
rect 1149 423 1152 429
rect 1140 417 1152 423
rect 1140 411 1143 417
rect 1149 411 1152 417
rect 1140 405 1152 411
rect 1140 399 1143 405
rect 1149 399 1152 405
rect 1140 396 1152 399
rect 1188 417 1200 432
rect 1188 411 1191 417
rect 1197 411 1200 417
rect 1188 405 1200 411
rect 1188 399 1191 405
rect 1197 399 1200 405
rect 1188 396 1200 399
rect 1236 429 1248 432
rect 1236 423 1239 429
rect 1245 423 1248 429
rect 1236 417 1248 423
rect 1236 411 1239 417
rect 1245 411 1248 417
rect 1236 405 1248 411
rect 1236 399 1239 405
rect 1245 399 1248 405
rect 1236 396 1248 399
rect 1284 417 1296 432
rect 1284 411 1287 417
rect 1293 411 1296 417
rect 1284 405 1296 411
rect 1284 399 1287 405
rect 1293 399 1296 405
rect 1284 396 1296 399
rect 1332 429 1344 432
rect 1332 423 1335 429
rect 1341 423 1344 429
rect 1332 417 1344 423
rect 1380 429 1392 432
rect 1380 423 1383 429
rect 1389 423 1392 429
rect 1332 411 1335 417
rect 1341 411 1344 417
rect 1332 405 1344 411
rect 1332 399 1335 405
rect 1341 399 1344 405
rect 1332 396 1344 399
rect 1356 417 1368 420
rect 1356 411 1359 417
rect 1365 411 1368 417
rect 1356 405 1368 411
rect 1356 399 1359 405
rect 1365 399 1368 405
rect 1356 396 1368 399
rect 1380 417 1392 423
rect 1428 429 1440 432
rect 1428 423 1431 429
rect 1437 423 1440 429
rect 1380 411 1383 417
rect 1389 411 1392 417
rect 1380 405 1392 411
rect 1380 399 1383 405
rect 1389 399 1392 405
rect 1380 396 1392 399
rect 1404 417 1416 420
rect 1404 411 1407 417
rect 1413 411 1416 417
rect 1404 405 1416 411
rect 1404 399 1407 405
rect 1413 399 1416 405
rect 1404 396 1416 399
rect 1428 417 1440 423
rect 1476 429 1488 432
rect 1476 423 1479 429
rect 1485 423 1488 429
rect 1428 411 1431 417
rect 1437 411 1440 417
rect 1428 405 1440 411
rect 1428 399 1431 405
rect 1437 399 1440 405
rect 1428 396 1440 399
rect 1452 417 1464 420
rect 1452 411 1455 417
rect 1461 411 1464 417
rect 1452 405 1464 411
rect 1452 399 1455 405
rect 1461 399 1464 405
rect 1452 396 1464 399
rect 1476 417 1488 423
rect 1524 429 1536 432
rect 1524 423 1527 429
rect 1533 423 1536 429
rect 1476 411 1479 417
rect 1485 411 1488 417
rect 1476 405 1488 411
rect 1476 399 1479 405
rect 1485 399 1488 405
rect 1476 396 1488 399
rect 1500 417 1512 420
rect 1500 411 1503 417
rect 1509 411 1512 417
rect 1500 405 1512 411
rect 1500 399 1503 405
rect 1509 399 1512 405
rect 1500 396 1512 399
rect 1524 417 1536 423
rect 1572 429 1584 432
rect 1572 423 1575 429
rect 1581 423 1584 429
rect 1524 411 1527 417
rect 1533 411 1536 417
rect 1524 405 1536 411
rect 1524 399 1527 405
rect 1533 399 1536 405
rect 1524 396 1536 399
rect 1548 417 1560 420
rect 1548 411 1551 417
rect 1557 411 1560 417
rect 1548 405 1560 411
rect 1548 399 1551 405
rect 1557 399 1560 405
rect 1548 384 1560 399
rect 1572 417 1584 423
rect 1572 411 1575 417
rect 1581 411 1584 417
rect 1572 405 1584 411
rect 1572 399 1575 405
rect 1581 399 1584 405
rect 1572 396 1584 399
rect 1596 429 1608 435
rect 1596 423 1599 429
rect 1605 423 1608 429
rect 1596 417 1608 423
rect 1596 411 1599 417
rect 1605 411 1608 417
rect 1596 405 1608 411
rect 1596 399 1599 405
rect 1605 399 1608 405
rect 1596 393 1608 399
rect 1596 387 1599 393
rect 1605 387 1608 393
rect -84 375 -81 381
rect -75 375 -72 381
rect -84 369 -72 375
rect -48 381 -12 384
rect -48 375 -45 381
rect -39 375 -33 381
rect -27 375 -21 381
rect -15 375 -12 381
rect -48 372 -12 375
rect 0 381 36 384
rect 0 375 3 381
rect 9 375 15 381
rect 21 375 27 381
rect 33 375 36 381
rect 0 372 36 375
rect 48 381 84 384
rect 48 375 51 381
rect 57 375 63 381
rect 69 375 75 381
rect 81 375 84 381
rect 48 372 84 375
rect 96 381 132 384
rect 96 375 99 381
rect 105 375 111 381
rect 117 375 123 381
rect 129 375 132 381
rect 96 372 132 375
rect 144 381 180 384
rect 144 375 147 381
rect 153 375 159 381
rect 165 375 171 381
rect 177 375 180 381
rect 144 372 180 375
rect 192 381 228 384
rect 192 375 195 381
rect 201 375 207 381
rect 213 375 219 381
rect 225 375 228 381
rect 192 372 228 375
rect 240 381 276 384
rect 240 375 243 381
rect 249 375 255 381
rect 261 375 267 381
rect 273 375 276 381
rect 240 372 276 375
rect 288 381 324 384
rect 288 375 291 381
rect 297 375 303 381
rect 309 375 315 381
rect 321 375 324 381
rect 288 372 324 375
rect 336 381 372 384
rect 336 375 339 381
rect 345 375 351 381
rect 357 375 363 381
rect 369 375 372 381
rect 336 372 372 375
rect 384 381 420 384
rect 384 375 387 381
rect 393 375 399 381
rect 405 375 411 381
rect 417 375 420 381
rect 384 372 420 375
rect 432 381 468 384
rect 432 375 435 381
rect 441 375 447 381
rect 453 375 459 381
rect 465 375 468 381
rect 432 372 468 375
rect 480 381 516 384
rect 480 375 483 381
rect 489 375 495 381
rect 501 375 507 381
rect 513 375 516 381
rect 480 372 516 375
rect 528 381 564 384
rect 528 375 531 381
rect 537 375 543 381
rect 549 375 555 381
rect 561 375 564 381
rect 528 372 564 375
rect 576 381 612 384
rect 576 375 579 381
rect 585 375 591 381
rect 597 375 603 381
rect 609 375 612 381
rect 576 372 612 375
rect 624 381 660 384
rect 624 375 627 381
rect 633 375 639 381
rect 645 375 651 381
rect 657 375 660 381
rect 624 372 660 375
rect 672 381 708 384
rect 672 375 675 381
rect 681 375 687 381
rect 693 375 699 381
rect 705 375 708 381
rect 672 372 708 375
rect 720 381 756 384
rect 720 375 723 381
rect 729 375 735 381
rect 741 375 747 381
rect 753 375 756 381
rect 720 372 756 375
rect 768 381 804 384
rect 768 375 771 381
rect 777 375 783 381
rect 789 375 795 381
rect 801 375 804 381
rect 768 372 804 375
rect 816 381 852 384
rect 816 375 819 381
rect 825 375 831 381
rect 837 375 843 381
rect 849 375 852 381
rect 816 372 852 375
rect 864 381 900 384
rect 864 375 867 381
rect 873 375 879 381
rect 885 375 891 381
rect 897 375 900 381
rect 864 372 900 375
rect 912 381 948 384
rect 912 375 915 381
rect 921 375 927 381
rect 933 375 939 381
rect 945 375 948 381
rect 912 372 948 375
rect 960 381 996 384
rect 960 375 963 381
rect 969 375 975 381
rect 981 375 987 381
rect 993 375 996 381
rect 960 372 996 375
rect 1008 381 1044 384
rect 1008 375 1011 381
rect 1017 375 1023 381
rect 1029 375 1035 381
rect 1041 375 1044 381
rect 1008 372 1044 375
rect 1056 381 1092 384
rect 1056 375 1059 381
rect 1065 375 1071 381
rect 1077 375 1083 381
rect 1089 375 1092 381
rect 1056 372 1092 375
rect 1104 381 1140 384
rect 1104 375 1107 381
rect 1113 375 1119 381
rect 1125 375 1131 381
rect 1137 375 1140 381
rect 1104 372 1140 375
rect 1152 381 1188 384
rect 1152 375 1155 381
rect 1161 375 1167 381
rect 1173 375 1179 381
rect 1185 375 1188 381
rect 1152 372 1188 375
rect 1200 381 1236 384
rect 1200 375 1203 381
rect 1209 375 1215 381
rect 1221 375 1227 381
rect 1233 375 1236 381
rect 1200 372 1236 375
rect 1248 381 1284 384
rect 1248 375 1251 381
rect 1257 375 1263 381
rect 1269 375 1275 381
rect 1281 375 1284 381
rect 1248 372 1284 375
rect 1296 381 1332 384
rect 1296 375 1299 381
rect 1305 375 1311 381
rect 1317 375 1323 381
rect 1329 375 1332 381
rect 1296 372 1332 375
rect 1344 381 1380 384
rect 1344 375 1347 381
rect 1353 375 1359 381
rect 1365 375 1371 381
rect 1377 375 1380 381
rect 1344 372 1380 375
rect 1392 381 1428 384
rect 1392 375 1395 381
rect 1401 375 1407 381
rect 1413 375 1419 381
rect 1425 375 1428 381
rect 1392 372 1428 375
rect 1440 381 1476 384
rect 1440 375 1443 381
rect 1449 375 1455 381
rect 1461 375 1467 381
rect 1473 375 1476 381
rect 1440 372 1476 375
rect 1488 381 1524 384
rect 1488 375 1491 381
rect 1497 375 1503 381
rect 1509 375 1515 381
rect 1521 375 1524 381
rect 1488 372 1524 375
rect 1536 381 1572 384
rect 1536 375 1539 381
rect 1545 375 1551 381
rect 1557 375 1563 381
rect 1569 375 1572 381
rect 1536 372 1572 375
rect 1596 381 1608 387
rect 1596 375 1599 381
rect 1605 375 1608 381
rect -84 363 -81 369
rect -75 363 -72 369
rect -84 360 -72 363
rect 1596 369 1608 375
rect 1596 363 1599 369
rect 1605 363 1608 369
rect 1596 360 1608 363
rect -84 357 1608 360
rect -84 351 -81 357
rect -75 351 -69 357
rect -63 351 -57 357
rect -51 351 -45 357
rect -39 351 -33 357
rect -27 351 -21 357
rect -15 351 -9 357
rect -3 351 3 357
rect 9 351 15 357
rect 21 351 27 357
rect 33 351 39 357
rect 45 351 51 357
rect 57 351 63 357
rect 69 351 75 357
rect 81 351 87 357
rect 93 351 99 357
rect 105 351 111 357
rect 117 351 123 357
rect 129 351 135 357
rect 141 351 147 357
rect 153 351 159 357
rect 165 351 171 357
rect 177 351 183 357
rect 189 351 195 357
rect 201 351 207 357
rect 213 351 219 357
rect 225 351 231 357
rect 237 351 243 357
rect 249 351 255 357
rect 261 351 267 357
rect 273 351 279 357
rect 285 351 291 357
rect 297 351 303 357
rect 309 351 315 357
rect 321 351 327 357
rect 333 351 339 357
rect 345 351 351 357
rect 357 351 363 357
rect 369 351 375 357
rect 381 351 387 357
rect 393 351 399 357
rect 405 351 411 357
rect 417 351 423 357
rect 429 351 435 357
rect 441 351 447 357
rect 453 351 459 357
rect 465 351 471 357
rect 477 351 483 357
rect 489 351 495 357
rect 501 351 507 357
rect 513 351 519 357
rect 525 351 531 357
rect 537 351 543 357
rect 549 351 555 357
rect 561 351 567 357
rect 573 351 579 357
rect 585 351 591 357
rect 597 351 603 357
rect 609 351 615 357
rect 621 351 627 357
rect 633 351 639 357
rect 645 351 651 357
rect 657 351 663 357
rect 669 351 675 357
rect 681 351 687 357
rect 693 351 699 357
rect 705 351 711 357
rect 717 351 723 357
rect 729 351 735 357
rect 741 351 747 357
rect 753 351 759 357
rect 765 351 771 357
rect 777 351 783 357
rect 789 351 795 357
rect 801 351 807 357
rect 813 351 819 357
rect 825 351 831 357
rect 837 351 843 357
rect 849 351 855 357
rect 861 351 867 357
rect 873 351 879 357
rect 885 351 891 357
rect 897 351 903 357
rect 909 351 915 357
rect 921 351 927 357
rect 933 351 939 357
rect 945 351 951 357
rect 957 351 963 357
rect 969 351 975 357
rect 981 351 987 357
rect 993 351 999 357
rect 1005 351 1011 357
rect 1017 351 1023 357
rect 1029 351 1035 357
rect 1041 351 1047 357
rect 1053 351 1059 357
rect 1065 351 1071 357
rect 1077 351 1083 357
rect 1089 351 1095 357
rect 1101 351 1107 357
rect 1113 351 1119 357
rect 1125 351 1131 357
rect 1137 351 1143 357
rect 1149 351 1155 357
rect 1161 351 1167 357
rect 1173 351 1179 357
rect 1185 351 1191 357
rect 1197 351 1203 357
rect 1209 351 1215 357
rect 1221 351 1227 357
rect 1233 351 1239 357
rect 1245 351 1251 357
rect 1257 351 1263 357
rect 1269 351 1275 357
rect 1281 351 1287 357
rect 1293 351 1299 357
rect 1305 351 1311 357
rect 1317 351 1323 357
rect 1329 351 1335 357
rect 1341 351 1347 357
rect 1353 351 1359 357
rect 1365 351 1371 357
rect 1377 351 1383 357
rect 1389 351 1395 357
rect 1401 351 1407 357
rect 1413 351 1419 357
rect 1425 351 1431 357
rect 1437 351 1443 357
rect 1449 351 1455 357
rect 1461 351 1467 357
rect 1473 351 1479 357
rect 1485 351 1491 357
rect 1497 351 1503 357
rect 1509 351 1515 357
rect 1521 351 1527 357
rect 1533 351 1539 357
rect 1545 351 1551 357
rect 1557 351 1563 357
rect 1569 351 1575 357
rect 1581 351 1587 357
rect 1593 351 1599 357
rect 1605 351 1608 357
rect -84 348 1608 351
rect 1620 453 1632 459
rect 1620 447 1623 453
rect 1629 447 1632 453
rect 1620 441 1632 447
rect 1620 435 1623 441
rect 1629 435 1632 441
rect 1620 429 1632 435
rect 1620 423 1623 429
rect 1629 423 1632 429
rect 1620 417 1632 423
rect 1620 411 1623 417
rect 1629 411 1632 417
rect 1620 405 1632 411
rect 1620 399 1623 405
rect 1629 399 1632 405
rect 1620 393 1632 399
rect 1620 387 1623 393
rect 1629 387 1632 393
rect 1620 381 1632 387
rect 1620 375 1623 381
rect 1629 375 1632 381
rect 1620 369 1632 375
rect 1620 363 1623 369
rect 1629 363 1632 369
rect 1620 357 1632 363
rect 1620 351 1623 357
rect 1629 351 1632 357
rect -108 339 -105 345
rect -99 339 -96 345
rect -108 336 -96 339
rect 1620 345 1632 351
rect 1620 339 1623 345
rect 1629 339 1632 345
rect 1620 336 1632 339
rect -108 333 1632 336
rect -108 327 -105 333
rect -99 327 -93 333
rect -87 327 -81 333
rect -75 327 -69 333
rect -63 327 -57 333
rect -51 327 -45 333
rect -39 327 -33 333
rect -27 327 -21 333
rect -15 327 -9 333
rect -3 327 3 333
rect 9 327 15 333
rect 21 327 27 333
rect 33 327 39 333
rect 45 327 51 333
rect 57 327 63 333
rect 69 327 75 333
rect 81 327 87 333
rect 93 327 99 333
rect 105 327 111 333
rect 117 327 123 333
rect 129 327 135 333
rect 141 327 147 333
rect 153 327 159 333
rect 165 327 171 333
rect 177 327 183 333
rect 189 327 195 333
rect 201 327 207 333
rect 213 327 219 333
rect 225 327 231 333
rect 237 327 243 333
rect 249 327 255 333
rect 261 327 267 333
rect 273 327 279 333
rect 285 327 291 333
rect 297 327 303 333
rect 309 327 315 333
rect 321 327 327 333
rect 333 327 339 333
rect 345 327 351 333
rect 357 327 363 333
rect 369 327 375 333
rect 381 327 387 333
rect 393 327 399 333
rect 405 327 411 333
rect 417 327 423 333
rect 429 327 435 333
rect 441 327 447 333
rect 453 327 459 333
rect 465 327 471 333
rect 477 327 483 333
rect 489 327 495 333
rect 501 327 507 333
rect 513 327 519 333
rect 525 327 531 333
rect 537 327 543 333
rect 549 327 555 333
rect 561 327 567 333
rect 573 327 579 333
rect 585 327 591 333
rect 597 327 603 333
rect 609 327 615 333
rect 621 327 627 333
rect 633 327 639 333
rect 645 327 651 333
rect 657 327 663 333
rect 669 327 675 333
rect 681 327 687 333
rect 693 327 699 333
rect 705 327 711 333
rect 717 327 723 333
rect 729 327 735 333
rect 741 327 747 333
rect 753 327 759 333
rect 765 327 771 333
rect 777 327 783 333
rect 789 327 795 333
rect 801 327 807 333
rect 813 327 819 333
rect 825 327 831 333
rect 837 327 843 333
rect 849 327 855 333
rect 861 327 867 333
rect 873 327 879 333
rect 885 327 891 333
rect 897 327 903 333
rect 909 327 915 333
rect 921 327 927 333
rect 933 327 939 333
rect 945 327 951 333
rect 957 327 963 333
rect 969 327 975 333
rect 981 327 987 333
rect 993 327 999 333
rect 1005 327 1011 333
rect 1017 327 1023 333
rect 1029 327 1035 333
rect 1041 327 1047 333
rect 1053 327 1059 333
rect 1065 327 1071 333
rect 1077 327 1083 333
rect 1089 327 1095 333
rect 1101 327 1107 333
rect 1113 327 1119 333
rect 1125 327 1131 333
rect 1137 327 1143 333
rect 1149 327 1155 333
rect 1161 327 1167 333
rect 1173 327 1179 333
rect 1185 327 1191 333
rect 1197 327 1203 333
rect 1209 327 1215 333
rect 1221 327 1227 333
rect 1233 327 1239 333
rect 1245 327 1251 333
rect 1257 327 1263 333
rect 1269 327 1275 333
rect 1281 327 1287 333
rect 1293 327 1299 333
rect 1305 327 1311 333
rect 1317 327 1323 333
rect 1329 327 1335 333
rect 1341 327 1347 333
rect 1353 327 1359 333
rect 1365 327 1371 333
rect 1377 327 1383 333
rect 1389 327 1395 333
rect 1401 327 1407 333
rect 1413 327 1419 333
rect 1425 327 1431 333
rect 1437 327 1443 333
rect 1449 327 1455 333
rect 1461 327 1467 333
rect 1473 327 1479 333
rect 1485 327 1491 333
rect 1497 327 1503 333
rect 1509 327 1515 333
rect 1521 327 1527 333
rect 1533 327 1539 333
rect 1545 327 1551 333
rect 1557 327 1563 333
rect 1569 327 1575 333
rect 1581 327 1587 333
rect 1593 327 1599 333
rect 1605 327 1611 333
rect 1617 327 1623 333
rect 1629 327 1632 333
rect -108 324 1632 327
rect -108 321 -96 324
rect -108 315 -105 321
rect -99 315 -96 321
rect -108 309 -96 315
rect -108 303 -105 309
rect -99 303 -96 309
rect -108 297 -96 303
rect -108 291 -105 297
rect -99 291 -96 297
rect -108 285 -96 291
rect -108 279 -105 285
rect -99 279 -96 285
rect -108 273 -96 279
rect -108 267 -105 273
rect -99 267 -96 273
rect -108 261 -96 267
rect -108 255 -105 261
rect -99 255 -96 261
rect -108 249 -96 255
rect -108 243 -105 249
rect -99 243 -96 249
rect -108 237 -96 243
rect -108 231 -105 237
rect -99 231 -96 237
rect -108 225 -96 231
rect -108 219 -105 225
rect -99 219 -96 225
rect -108 213 -96 219
rect -108 207 -105 213
rect -99 207 -96 213
rect -108 201 -96 207
rect -108 195 -105 201
rect -99 195 -96 201
rect -108 189 -96 195
rect -108 183 -105 189
rect -99 183 -96 189
rect -108 177 -96 183
rect -108 171 -105 177
rect -99 171 -96 177
rect -108 165 -96 171
rect -108 159 -105 165
rect -99 159 -96 165
rect -108 153 -96 159
rect -108 147 -105 153
rect -99 147 -96 153
rect -108 141 -96 147
rect -108 135 -105 141
rect -99 135 -96 141
rect -108 129 -96 135
rect -108 123 -105 129
rect -99 123 -96 129
rect -108 117 -96 123
rect -108 111 -105 117
rect -99 111 -96 117
rect -108 105 -96 111
rect -108 99 -105 105
rect -99 99 -96 105
rect -108 96 -96 99
rect 1620 321 1632 324
rect 1620 315 1623 321
rect 1629 315 1632 321
rect 1620 309 1632 315
rect 1620 303 1623 309
rect 1629 303 1632 309
rect 1620 297 1632 303
rect 1620 291 1623 297
rect 1629 291 1632 297
rect 1620 285 1632 291
rect 1620 279 1623 285
rect 1629 279 1632 285
rect 1620 273 1632 279
rect 1620 267 1623 273
rect 1629 267 1632 273
rect 1620 261 1632 267
rect 1620 255 1623 261
rect 1629 255 1632 261
rect 1620 249 1632 255
rect 1620 243 1623 249
rect 1629 243 1632 249
rect 1620 237 1632 243
rect 1620 231 1623 237
rect 1629 231 1632 237
rect 1620 225 1632 231
rect 1620 219 1623 225
rect 1629 219 1632 225
rect 1620 213 1632 219
rect 1620 207 1623 213
rect 1629 207 1632 213
rect 1620 201 1632 207
rect 1620 195 1623 201
rect 1629 195 1632 201
rect 1620 189 1632 195
rect 1620 183 1623 189
rect 1629 183 1632 189
rect 1620 177 1632 183
rect 1620 171 1623 177
rect 1629 171 1632 177
rect 1620 165 1632 171
rect 1620 159 1623 165
rect 1629 159 1632 165
rect 1620 153 1632 159
rect 1620 147 1623 153
rect 1629 147 1632 153
rect 1620 141 1632 147
rect 1620 135 1623 141
rect 1629 135 1632 141
rect 1620 129 1632 135
rect 1620 123 1623 129
rect 1629 123 1632 129
rect 1620 117 1632 123
rect 1620 111 1623 117
rect 1629 111 1632 117
rect 1620 105 1632 111
rect 1620 99 1623 105
rect 1629 99 1632 105
rect 1620 96 1632 99
rect -108 93 1632 96
rect -108 87 -105 93
rect -99 87 -93 93
rect -87 87 -81 93
rect -75 87 -69 93
rect -63 87 -57 93
rect -51 87 -45 93
rect -39 87 -33 93
rect -27 87 -21 93
rect -15 87 -9 93
rect -3 87 3 93
rect 9 87 15 93
rect 21 87 27 93
rect 33 87 39 93
rect 45 87 51 93
rect 57 87 63 93
rect 69 87 75 93
rect 81 87 87 93
rect 93 87 99 93
rect 105 87 111 93
rect 117 87 123 93
rect 129 87 135 93
rect 141 87 147 93
rect 153 87 159 93
rect 165 87 171 93
rect 177 87 183 93
rect 189 87 195 93
rect 201 87 207 93
rect 213 87 219 93
rect 225 87 231 93
rect 237 87 243 93
rect 249 87 255 93
rect 261 87 267 93
rect 273 87 279 93
rect 285 87 291 93
rect 297 87 303 93
rect 309 87 315 93
rect 321 87 327 93
rect 333 87 339 93
rect 345 87 351 93
rect 357 87 363 93
rect 369 87 375 93
rect 381 87 387 93
rect 393 87 399 93
rect 405 87 411 93
rect 417 87 423 93
rect 429 87 435 93
rect 441 87 447 93
rect 453 87 459 93
rect 465 87 471 93
rect 477 87 483 93
rect 489 87 495 93
rect 501 87 507 93
rect 513 87 519 93
rect 525 87 531 93
rect 537 87 543 93
rect 549 87 555 93
rect 561 87 567 93
rect 573 87 579 93
rect 585 87 591 93
rect 597 87 603 93
rect 609 87 615 93
rect 621 87 627 93
rect 633 87 639 93
rect 645 87 651 93
rect 657 87 663 93
rect 669 87 675 93
rect 681 87 687 93
rect 693 87 699 93
rect 705 87 711 93
rect 717 87 723 93
rect 729 87 735 93
rect 741 87 747 93
rect 753 87 759 93
rect 765 87 771 93
rect 777 87 783 93
rect 789 87 795 93
rect 801 87 807 93
rect 813 87 819 93
rect 825 87 831 93
rect 837 87 843 93
rect 849 87 855 93
rect 861 87 867 93
rect 873 87 879 93
rect 885 87 891 93
rect 897 87 903 93
rect 909 87 915 93
rect 921 87 927 93
rect 933 87 939 93
rect 945 87 951 93
rect 957 87 963 93
rect 969 87 975 93
rect 981 87 987 93
rect 993 87 999 93
rect 1005 87 1011 93
rect 1017 87 1023 93
rect 1029 87 1035 93
rect 1041 87 1047 93
rect 1053 87 1059 93
rect 1065 87 1071 93
rect 1077 87 1083 93
rect 1089 87 1095 93
rect 1101 87 1107 93
rect 1113 87 1119 93
rect 1125 87 1131 93
rect 1137 87 1143 93
rect 1149 87 1155 93
rect 1161 87 1167 93
rect 1173 87 1179 93
rect 1185 87 1191 93
rect 1197 87 1203 93
rect 1209 87 1215 93
rect 1221 87 1227 93
rect 1233 87 1239 93
rect 1245 87 1251 93
rect 1257 87 1263 93
rect 1269 87 1275 93
rect 1281 87 1287 93
rect 1293 87 1299 93
rect 1305 87 1311 93
rect 1317 87 1323 93
rect 1329 87 1335 93
rect 1341 87 1347 93
rect 1353 87 1359 93
rect 1365 87 1371 93
rect 1377 87 1383 93
rect 1389 87 1395 93
rect 1401 87 1407 93
rect 1413 87 1419 93
rect 1425 87 1431 93
rect 1437 87 1443 93
rect 1449 87 1455 93
rect 1461 87 1467 93
rect 1473 87 1479 93
rect 1485 87 1491 93
rect 1497 87 1503 93
rect 1509 87 1515 93
rect 1521 87 1527 93
rect 1533 87 1539 93
rect 1545 87 1551 93
rect 1557 87 1563 93
rect 1569 87 1575 93
rect 1581 87 1587 93
rect 1593 87 1599 93
rect 1605 87 1611 93
rect 1617 87 1623 93
rect 1629 87 1632 93
rect -108 84 1632 87
rect -108 81 -96 84
rect -108 75 -105 81
rect -99 75 -96 81
rect -108 69 -96 75
rect 1620 81 1632 84
rect 1620 75 1623 81
rect 1629 75 1632 81
rect -108 63 -105 69
rect -99 63 -96 69
rect -108 57 -96 63
rect -48 69 -12 72
rect -48 63 -45 69
rect -39 63 -33 69
rect -27 63 -21 69
rect -15 63 -12 69
rect -48 60 -12 63
rect 0 69 36 72
rect 0 63 3 69
rect 9 63 15 69
rect 21 63 27 69
rect 33 63 36 69
rect 0 60 36 63
rect 48 69 84 72
rect 48 63 51 69
rect 57 63 63 69
rect 69 63 75 69
rect 81 63 84 69
rect 48 60 84 63
rect 96 69 132 72
rect 96 63 99 69
rect 105 63 111 69
rect 117 63 123 69
rect 129 63 132 69
rect 96 60 132 63
rect 144 69 180 72
rect 144 63 147 69
rect 153 63 159 69
rect 165 63 171 69
rect 177 63 180 69
rect 144 60 180 63
rect 192 69 228 72
rect 192 63 195 69
rect 201 63 207 69
rect 213 63 219 69
rect 225 63 228 69
rect 192 60 228 63
rect 240 69 276 72
rect 240 63 243 69
rect 249 63 255 69
rect 261 63 267 69
rect 273 63 276 69
rect 240 60 276 63
rect 288 69 324 72
rect 288 63 291 69
rect 297 63 303 69
rect 309 63 315 69
rect 321 63 324 69
rect 288 60 324 63
rect 336 69 372 72
rect 336 63 339 69
rect 345 63 351 69
rect 357 63 363 69
rect 369 63 372 69
rect 336 60 372 63
rect 384 69 420 72
rect 384 63 387 69
rect 393 63 399 69
rect 405 63 411 69
rect 417 63 420 69
rect 384 60 420 63
rect 432 69 468 72
rect 432 63 435 69
rect 441 63 447 69
rect 453 63 459 69
rect 465 63 468 69
rect 432 60 468 63
rect 480 69 516 72
rect 480 63 483 69
rect 489 63 495 69
rect 501 63 507 69
rect 513 63 516 69
rect 480 60 516 63
rect 528 69 564 72
rect 528 63 531 69
rect 537 63 543 69
rect 549 63 555 69
rect 561 63 564 69
rect 528 60 564 63
rect 576 69 612 72
rect 576 63 579 69
rect 585 63 591 69
rect 597 63 603 69
rect 609 63 612 69
rect 576 60 612 63
rect 624 69 660 72
rect 624 63 627 69
rect 633 63 639 69
rect 645 63 651 69
rect 657 63 660 69
rect 624 60 660 63
rect 672 69 708 72
rect 672 63 675 69
rect 681 63 687 69
rect 693 63 699 69
rect 705 63 708 69
rect 672 60 708 63
rect 720 69 756 72
rect 720 63 723 69
rect 729 63 735 69
rect 741 63 747 69
rect 753 63 756 69
rect 720 60 756 63
rect 768 69 804 72
rect 768 63 771 69
rect 777 63 783 69
rect 789 63 795 69
rect 801 63 804 69
rect 768 60 804 63
rect 816 69 852 72
rect 816 63 819 69
rect 825 63 831 69
rect 837 63 843 69
rect 849 63 852 69
rect 816 60 852 63
rect 864 69 900 72
rect 864 63 867 69
rect 873 63 879 69
rect 885 63 891 69
rect 897 63 900 69
rect 864 60 900 63
rect 912 69 948 72
rect 912 63 915 69
rect 921 63 927 69
rect 933 63 939 69
rect 945 63 948 69
rect 912 60 948 63
rect 960 69 996 72
rect 960 63 963 69
rect 969 63 975 69
rect 981 63 987 69
rect 993 63 996 69
rect 960 60 996 63
rect 1008 69 1044 72
rect 1008 63 1011 69
rect 1017 63 1023 69
rect 1029 63 1035 69
rect 1041 63 1044 69
rect 1008 60 1044 63
rect 1056 69 1092 72
rect 1056 63 1059 69
rect 1065 63 1071 69
rect 1077 63 1083 69
rect 1089 63 1092 69
rect 1056 60 1092 63
rect 1104 69 1140 72
rect 1104 63 1107 69
rect 1113 63 1119 69
rect 1125 63 1131 69
rect 1137 63 1140 69
rect 1104 60 1140 63
rect 1152 69 1188 72
rect 1152 63 1155 69
rect 1161 63 1167 69
rect 1173 63 1179 69
rect 1185 63 1188 69
rect 1152 60 1188 63
rect 1200 69 1236 72
rect 1200 63 1203 69
rect 1209 63 1215 69
rect 1221 63 1227 69
rect 1233 63 1236 69
rect 1200 60 1236 63
rect 1248 69 1284 72
rect 1248 63 1251 69
rect 1257 63 1263 69
rect 1269 63 1275 69
rect 1281 63 1284 69
rect 1248 60 1284 63
rect 1296 69 1332 72
rect 1296 63 1299 69
rect 1305 63 1311 69
rect 1317 63 1323 69
rect 1329 63 1332 69
rect 1296 60 1332 63
rect 1344 69 1380 72
rect 1344 63 1347 69
rect 1353 63 1359 69
rect 1365 63 1371 69
rect 1377 63 1380 69
rect 1344 60 1380 63
rect 1392 69 1428 72
rect 1392 63 1395 69
rect 1401 63 1407 69
rect 1413 63 1419 69
rect 1425 63 1428 69
rect 1392 60 1428 63
rect 1440 69 1476 72
rect 1440 63 1443 69
rect 1449 63 1455 69
rect 1461 63 1467 69
rect 1473 63 1476 69
rect 1440 60 1476 63
rect 1488 69 1524 72
rect 1488 63 1491 69
rect 1497 63 1503 69
rect 1509 63 1515 69
rect 1521 63 1524 69
rect 1488 60 1524 63
rect 1536 69 1572 72
rect 1536 63 1539 69
rect 1545 63 1551 69
rect 1557 63 1563 69
rect 1569 63 1572 69
rect 1536 60 1572 63
rect 1620 69 1632 75
rect 1620 63 1623 69
rect 1629 63 1632 69
rect -108 51 -105 57
rect -99 51 -96 57
rect -108 45 -96 51
rect -108 39 -105 45
rect -99 39 -96 45
rect -108 33 -96 39
rect -108 27 -105 33
rect -99 27 -96 33
rect -108 21 -96 27
rect -108 15 -105 21
rect -99 15 -96 21
rect -108 9 -96 15
rect -60 45 -48 48
rect -60 39 -57 45
rect -51 39 -48 45
rect -60 33 -48 39
rect -60 27 -57 33
rect -51 27 -48 33
rect -60 21 -48 27
rect -60 15 -57 21
rect -51 15 -48 21
rect -60 12 -48 15
rect -36 45 -24 60
rect -36 39 -33 45
rect -27 39 -24 45
rect -36 33 -24 39
rect -36 27 -33 33
rect -27 27 -24 33
rect -36 21 -24 27
rect -36 15 -33 21
rect -27 15 -24 21
rect -36 12 -24 15
rect -12 45 0 48
rect -12 39 -9 45
rect -3 39 0 45
rect -12 33 0 39
rect -12 27 -9 33
rect -3 27 0 33
rect -12 21 0 27
rect -12 15 -9 21
rect -3 15 0 21
rect -12 12 0 15
rect 36 45 48 48
rect 36 39 39 45
rect 45 39 48 45
rect 36 33 48 39
rect 36 27 39 33
rect 45 27 48 33
rect 36 21 48 27
rect 36 15 39 21
rect 45 15 48 21
rect 36 12 48 15
rect 84 45 96 48
rect 84 39 87 45
rect 93 39 96 45
rect 84 33 96 39
rect 84 27 87 33
rect 93 27 96 33
rect 84 21 96 27
rect 84 15 87 21
rect 93 15 96 21
rect 84 12 96 15
rect 132 45 144 48
rect 132 39 135 45
rect 141 39 144 45
rect 132 33 144 39
rect 132 27 135 33
rect 141 27 144 33
rect 132 21 144 27
rect 132 15 135 21
rect 141 15 144 21
rect 132 12 144 15
rect 180 45 192 48
rect 180 39 183 45
rect 189 39 192 45
rect 180 33 192 39
rect 180 27 183 33
rect 189 27 192 33
rect 180 21 192 27
rect 180 15 183 21
rect 189 15 192 21
rect 180 12 192 15
rect 276 45 288 48
rect 276 39 279 45
rect 285 39 288 45
rect 276 33 288 39
rect 276 27 279 33
rect 285 27 288 33
rect 276 21 288 27
rect 276 15 279 21
rect 285 15 288 21
rect 276 12 288 15
rect 372 45 384 48
rect 372 39 375 45
rect 381 39 384 45
rect 372 33 384 39
rect 372 27 375 33
rect 381 27 384 33
rect 372 21 384 27
rect 372 15 375 21
rect 381 15 384 21
rect 372 12 384 15
rect 468 45 480 48
rect 468 39 471 45
rect 477 39 480 45
rect 468 33 480 39
rect 468 27 471 33
rect 477 27 480 33
rect 468 21 480 27
rect 468 15 471 21
rect 477 15 480 21
rect 468 12 480 15
rect 564 45 576 48
rect 564 39 567 45
rect 573 39 576 45
rect 564 33 576 39
rect 564 27 567 33
rect 573 27 576 33
rect 564 21 576 27
rect 564 15 567 21
rect 573 15 576 21
rect 564 12 576 15
rect 612 45 624 48
rect 612 39 615 45
rect 621 39 624 45
rect 612 33 624 39
rect 612 27 615 33
rect 621 27 624 33
rect 612 21 624 27
rect 612 15 615 21
rect 621 15 624 21
rect 612 12 624 15
rect 660 45 672 48
rect 660 39 663 45
rect 669 39 672 45
rect 660 33 672 39
rect 660 27 663 33
rect 669 27 672 33
rect 660 21 672 27
rect 660 15 663 21
rect 669 15 672 21
rect 660 12 672 15
rect 708 45 720 48
rect 708 39 711 45
rect 717 39 720 45
rect 708 33 720 39
rect 708 27 711 33
rect 717 27 720 33
rect 708 21 720 27
rect 708 15 711 21
rect 717 15 720 21
rect 708 12 720 15
rect 756 45 768 48
rect 756 39 759 45
rect 765 39 768 45
rect 756 33 768 39
rect 756 27 759 33
rect 765 27 768 33
rect 756 21 768 27
rect 756 15 759 21
rect 765 15 768 21
rect 756 12 768 15
rect 804 45 816 48
rect 804 39 807 45
rect 813 39 816 45
rect 804 33 816 39
rect 804 27 807 33
rect 813 27 816 33
rect 804 21 816 27
rect 804 15 807 21
rect 813 15 816 21
rect 804 12 816 15
rect 852 45 864 48
rect 852 39 855 45
rect 861 39 864 45
rect 852 33 864 39
rect 852 27 855 33
rect 861 27 864 33
rect 852 21 864 27
rect 852 15 855 21
rect 861 15 864 21
rect 852 12 864 15
rect 900 45 912 48
rect 900 39 903 45
rect 909 39 912 45
rect 900 33 912 39
rect 900 27 903 33
rect 909 27 912 33
rect 900 21 912 27
rect 900 15 903 21
rect 909 15 912 21
rect 900 12 912 15
rect 948 45 960 48
rect 948 39 951 45
rect 957 39 960 45
rect 948 33 960 39
rect 948 27 951 33
rect 957 27 960 33
rect 948 21 960 27
rect 948 15 951 21
rect 957 15 960 21
rect 948 12 960 15
rect 1044 45 1056 48
rect 1044 39 1047 45
rect 1053 39 1056 45
rect 1044 33 1056 39
rect 1044 27 1047 33
rect 1053 27 1056 33
rect 1044 21 1056 27
rect 1044 15 1047 21
rect 1053 15 1056 21
rect 1044 12 1056 15
rect 1140 45 1152 48
rect 1140 39 1143 45
rect 1149 39 1152 45
rect 1140 33 1152 39
rect 1140 27 1143 33
rect 1149 27 1152 33
rect 1140 21 1152 27
rect 1140 15 1143 21
rect 1149 15 1152 21
rect 1140 12 1152 15
rect 1236 45 1248 48
rect 1236 39 1239 45
rect 1245 39 1248 45
rect 1236 33 1248 39
rect 1236 27 1239 33
rect 1245 27 1248 33
rect 1236 21 1248 27
rect 1236 15 1239 21
rect 1245 15 1248 21
rect 1236 12 1248 15
rect 1332 45 1344 48
rect 1332 39 1335 45
rect 1341 39 1344 45
rect 1332 33 1344 39
rect 1332 27 1335 33
rect 1341 27 1344 33
rect 1332 21 1344 27
rect 1332 15 1335 21
rect 1341 15 1344 21
rect 1332 12 1344 15
rect 1380 45 1392 48
rect 1380 39 1383 45
rect 1389 39 1392 45
rect 1380 33 1392 39
rect 1380 27 1383 33
rect 1389 27 1392 33
rect 1380 21 1392 27
rect 1380 15 1383 21
rect 1389 15 1392 21
rect 1380 12 1392 15
rect 1428 45 1440 48
rect 1428 39 1431 45
rect 1437 39 1440 45
rect 1428 33 1440 39
rect 1428 27 1431 33
rect 1437 27 1440 33
rect 1428 21 1440 27
rect 1428 15 1431 21
rect 1437 15 1440 21
rect 1428 12 1440 15
rect 1476 45 1488 48
rect 1476 39 1479 45
rect 1485 39 1488 45
rect 1476 33 1488 39
rect 1476 27 1479 33
rect 1485 27 1488 33
rect 1476 21 1488 27
rect 1476 15 1479 21
rect 1485 15 1488 21
rect 1476 12 1488 15
rect 1524 45 1536 48
rect 1524 39 1527 45
rect 1533 39 1536 45
rect 1524 33 1536 39
rect 1524 27 1527 33
rect 1533 27 1536 33
rect 1524 21 1536 27
rect 1524 15 1527 21
rect 1533 15 1536 21
rect 1524 12 1536 15
rect 1548 45 1560 60
rect 1620 57 1632 63
rect 1620 51 1623 57
rect 1629 51 1632 57
rect 1548 39 1551 45
rect 1557 39 1560 45
rect 1548 33 1560 39
rect 1548 27 1551 33
rect 1557 27 1560 33
rect 1548 21 1560 27
rect 1548 15 1551 21
rect 1557 15 1560 21
rect 1548 12 1560 15
rect 1572 45 1584 48
rect 1572 39 1575 45
rect 1581 39 1584 45
rect 1572 33 1584 39
rect 1572 27 1575 33
rect 1581 27 1584 33
rect 1572 21 1584 27
rect 1572 15 1575 21
rect 1581 15 1584 21
rect 1572 12 1584 15
rect 1620 45 1632 51
rect 1620 39 1623 45
rect 1629 39 1632 45
rect 1620 33 1632 39
rect 1620 27 1623 33
rect 1629 27 1632 33
rect 1620 21 1632 27
rect 1620 15 1623 21
rect 1629 15 1632 21
rect -108 3 -105 9
rect -99 3 -96 9
rect -108 0 -96 3
rect 1620 9 1632 15
rect 1620 3 1623 9
rect 1629 3 1632 9
rect 1620 0 1632 3
rect -108 -3 1632 0
rect -108 -9 -105 -3
rect -99 -9 -93 -3
rect -87 -9 -81 -3
rect -75 -9 -69 -3
rect -63 -9 -57 -3
rect -51 -9 -45 -3
rect -39 -9 -33 -3
rect -27 -9 -21 -3
rect -15 -9 -9 -3
rect -3 -9 3 -3
rect 9 -9 15 -3
rect 21 -9 27 -3
rect 33 -9 39 -3
rect 45 -9 51 -3
rect 57 -9 63 -3
rect 69 -9 75 -3
rect 81 -9 87 -3
rect 93 -9 99 -3
rect 105 -9 111 -3
rect 117 -9 123 -3
rect 129 -9 135 -3
rect 141 -9 147 -3
rect 153 -9 159 -3
rect 165 -9 171 -3
rect 177 -9 183 -3
rect 189 -9 195 -3
rect 201 -9 207 -3
rect 213 -9 219 -3
rect 225 -9 231 -3
rect 237 -9 243 -3
rect 249 -9 255 -3
rect 261 -9 267 -3
rect 273 -9 279 -3
rect 285 -9 291 -3
rect 297 -9 303 -3
rect 309 -9 315 -3
rect 321 -9 327 -3
rect 333 -9 339 -3
rect 345 -9 351 -3
rect 357 -9 363 -3
rect 369 -9 375 -3
rect 381 -9 387 -3
rect 393 -9 399 -3
rect 405 -9 411 -3
rect 417 -9 423 -3
rect 429 -9 435 -3
rect 441 -9 447 -3
rect 453 -9 459 -3
rect 465 -9 471 -3
rect 477 -9 483 -3
rect 489 -9 495 -3
rect 501 -9 507 -3
rect 513 -9 519 -3
rect 525 -9 531 -3
rect 537 -9 543 -3
rect 549 -9 555 -3
rect 561 -9 567 -3
rect 573 -9 579 -3
rect 585 -9 591 -3
rect 597 -9 603 -3
rect 609 -9 615 -3
rect 621 -9 627 -3
rect 633 -9 639 -3
rect 645 -9 651 -3
rect 657 -9 663 -3
rect 669 -9 675 -3
rect 681 -9 687 -3
rect 693 -9 699 -3
rect 705 -9 711 -3
rect 717 -9 723 -3
rect 729 -9 735 -3
rect 741 -9 747 -3
rect 753 -9 759 -3
rect 765 -9 771 -3
rect 777 -9 783 -3
rect 789 -9 795 -3
rect 801 -9 807 -3
rect 813 -9 819 -3
rect 825 -9 831 -3
rect 837 -9 843 -3
rect 849 -9 855 -3
rect 861 -9 867 -3
rect 873 -9 879 -3
rect 885 -9 891 -3
rect 897 -9 903 -3
rect 909 -9 915 -3
rect 921 -9 927 -3
rect 933 -9 939 -3
rect 945 -9 951 -3
rect 957 -9 963 -3
rect 969 -9 975 -3
rect 981 -9 987 -3
rect 993 -9 999 -3
rect 1005 -9 1011 -3
rect 1017 -9 1023 -3
rect 1029 -9 1035 -3
rect 1041 -9 1047 -3
rect 1053 -9 1059 -3
rect 1065 -9 1071 -3
rect 1077 -9 1083 -3
rect 1089 -9 1095 -3
rect 1101 -9 1107 -3
rect 1113 -9 1119 -3
rect 1125 -9 1131 -3
rect 1137 -9 1143 -3
rect 1149 -9 1155 -3
rect 1161 -9 1167 -3
rect 1173 -9 1179 -3
rect 1185 -9 1191 -3
rect 1197 -9 1203 -3
rect 1209 -9 1215 -3
rect 1221 -9 1227 -3
rect 1233 -9 1239 -3
rect 1245 -9 1251 -3
rect 1257 -9 1263 -3
rect 1269 -9 1275 -3
rect 1281 -9 1287 -3
rect 1293 -9 1299 -3
rect 1305 -9 1311 -3
rect 1317 -9 1323 -3
rect 1329 -9 1335 -3
rect 1341 -9 1347 -3
rect 1353 -9 1359 -3
rect 1365 -9 1371 -3
rect 1377 -9 1383 -3
rect 1389 -9 1395 -3
rect 1401 -9 1407 -3
rect 1413 -9 1419 -3
rect 1425 -9 1431 -3
rect 1437 -9 1443 -3
rect 1449 -9 1455 -3
rect 1461 -9 1467 -3
rect 1473 -9 1479 -3
rect 1485 -9 1491 -3
rect 1497 -9 1503 -3
rect 1509 -9 1515 -3
rect 1521 -9 1527 -3
rect 1533 -9 1539 -3
rect 1545 -9 1551 -3
rect 1557 -9 1563 -3
rect 1569 -9 1575 -3
rect 1581 -9 1587 -3
rect 1593 -9 1599 -3
rect 1605 -9 1611 -3
rect 1617 -9 1623 -3
rect 1629 -9 1632 -3
rect -108 -12 1632 -9
rect -108 -15 -96 -12
rect -108 -21 -105 -15
rect -99 -21 -96 -15
rect -108 -27 -96 -21
rect -108 -33 -105 -27
rect -99 -33 -96 -27
rect -108 -39 -96 -33
rect -108 -45 -105 -39
rect -99 -45 -96 -39
rect -108 -51 -96 -45
rect -108 -57 -105 -51
rect -99 -57 -96 -51
rect -108 -63 -96 -57
rect -108 -69 -105 -63
rect -99 -69 -96 -63
rect -108 -75 -96 -69
rect -108 -81 -105 -75
rect -99 -81 -96 -75
rect -108 -87 -96 -81
rect -108 -93 -105 -87
rect -99 -93 -96 -87
rect -108 -99 -96 -93
rect -108 -105 -105 -99
rect -99 -105 -96 -99
rect -108 -111 -96 -105
rect -108 -117 -105 -111
rect -99 -117 -96 -111
rect -108 -123 -96 -117
rect -108 -129 -105 -123
rect -99 -129 -96 -123
rect -108 -135 -96 -129
rect -108 -141 -105 -135
rect -99 -141 -96 -135
rect -108 -147 -96 -141
rect -108 -153 -105 -147
rect -99 -153 -96 -147
rect -108 -159 -96 -153
rect -108 -165 -105 -159
rect -99 -165 -96 -159
rect -108 -171 -96 -165
rect -108 -177 -105 -171
rect -99 -177 -96 -171
rect -108 -183 -96 -177
rect -108 -189 -105 -183
rect -99 -189 -96 -183
rect -108 -192 -96 -189
rect 1620 -15 1632 -12
rect 1620 -21 1623 -15
rect 1629 -21 1632 -15
rect 1620 -27 1632 -21
rect 1620 -33 1623 -27
rect 1629 -33 1632 -27
rect 1620 -39 1632 -33
rect 1620 -45 1623 -39
rect 1629 -45 1632 -39
rect 1620 -51 1632 -45
rect 1620 -57 1623 -51
rect 1629 -57 1632 -51
rect 1620 -63 1632 -57
rect 1620 -69 1623 -63
rect 1629 -69 1632 -63
rect 1620 -75 1632 -69
rect 1620 -81 1623 -75
rect 1629 -81 1632 -75
rect 1620 -87 1632 -81
rect 1620 -93 1623 -87
rect 1629 -93 1632 -87
rect 1620 -99 1632 -93
rect 1620 -105 1623 -99
rect 1629 -105 1632 -99
rect 1620 -111 1632 -105
rect 1620 -117 1623 -111
rect 1629 -117 1632 -111
rect 1620 -123 1632 -117
rect 1620 -129 1623 -123
rect 1629 -129 1632 -123
rect 1620 -135 1632 -129
rect 1620 -141 1623 -135
rect 1629 -141 1632 -135
rect 1620 -147 1632 -141
rect 1620 -153 1623 -147
rect 1629 -153 1632 -147
rect 1620 -159 1632 -153
rect 1620 -165 1623 -159
rect 1629 -165 1632 -159
rect 1620 -171 1632 -165
rect 1620 -177 1623 -171
rect 1629 -177 1632 -171
rect 1620 -183 1632 -177
rect 1620 -189 1623 -183
rect 1629 -189 1632 -183
rect 1620 -192 1632 -189
rect -108 -195 1632 -192
rect -108 -201 -105 -195
rect -99 -201 -93 -195
rect -87 -201 -81 -195
rect -75 -201 -69 -195
rect -63 -201 -57 -195
rect -51 -201 -45 -195
rect -39 -201 -33 -195
rect -27 -201 -21 -195
rect -15 -201 -9 -195
rect -3 -201 3 -195
rect 9 -201 15 -195
rect 21 -201 27 -195
rect 33 -201 39 -195
rect 45 -201 51 -195
rect 57 -201 63 -195
rect 69 -201 75 -195
rect 81 -201 87 -195
rect 93 -201 99 -195
rect 105 -201 111 -195
rect 117 -201 123 -195
rect 129 -201 135 -195
rect 141 -201 147 -195
rect 153 -201 159 -195
rect 165 -201 171 -195
rect 177 -201 183 -195
rect 189 -201 195 -195
rect 201 -201 207 -195
rect 213 -201 219 -195
rect 225 -201 231 -195
rect 237 -201 243 -195
rect 249 -201 255 -195
rect 261 -201 267 -195
rect 273 -201 279 -195
rect 285 -201 291 -195
rect 297 -201 303 -195
rect 309 -201 315 -195
rect 321 -201 327 -195
rect 333 -201 339 -195
rect 345 -201 351 -195
rect 357 -201 363 -195
rect 369 -201 375 -195
rect 381 -201 387 -195
rect 393 -201 399 -195
rect 405 -201 411 -195
rect 417 -201 423 -195
rect 429 -201 435 -195
rect 441 -201 447 -195
rect 453 -201 459 -195
rect 465 -201 471 -195
rect 477 -201 483 -195
rect 489 -201 495 -195
rect 501 -201 507 -195
rect 513 -201 519 -195
rect 525 -201 531 -195
rect 537 -201 543 -195
rect 549 -201 555 -195
rect 561 -201 567 -195
rect 573 -201 579 -195
rect 585 -201 591 -195
rect 597 -201 603 -195
rect 609 -201 615 -195
rect 621 -201 627 -195
rect 633 -201 639 -195
rect 645 -201 651 -195
rect 657 -201 663 -195
rect 669 -201 675 -195
rect 681 -201 687 -195
rect 693 -201 699 -195
rect 705 -201 711 -195
rect 717 -201 723 -195
rect 729 -201 735 -195
rect 741 -201 747 -195
rect 753 -201 759 -195
rect 765 -201 771 -195
rect 777 -201 783 -195
rect 789 -201 795 -195
rect 801 -201 807 -195
rect 813 -201 819 -195
rect 825 -201 831 -195
rect 837 -201 843 -195
rect 849 -201 855 -195
rect 861 -201 867 -195
rect 873 -201 879 -195
rect 885 -201 891 -195
rect 897 -201 903 -195
rect 909 -201 915 -195
rect 921 -201 927 -195
rect 933 -201 939 -195
rect 945 -201 951 -195
rect 957 -201 963 -195
rect 969 -201 975 -195
rect 981 -201 987 -195
rect 993 -201 999 -195
rect 1005 -201 1011 -195
rect 1017 -201 1023 -195
rect 1029 -201 1035 -195
rect 1041 -201 1047 -195
rect 1053 -201 1059 -195
rect 1065 -201 1071 -195
rect 1077 -201 1083 -195
rect 1089 -201 1095 -195
rect 1101 -201 1107 -195
rect 1113 -201 1119 -195
rect 1125 -201 1131 -195
rect 1137 -201 1143 -195
rect 1149 -201 1155 -195
rect 1161 -201 1167 -195
rect 1173 -201 1179 -195
rect 1185 -201 1191 -195
rect 1197 -201 1203 -195
rect 1209 -201 1215 -195
rect 1221 -201 1227 -195
rect 1233 -201 1239 -195
rect 1245 -201 1251 -195
rect 1257 -201 1263 -195
rect 1269 -201 1275 -195
rect 1281 -201 1287 -195
rect 1293 -201 1299 -195
rect 1305 -201 1311 -195
rect 1317 -201 1323 -195
rect 1329 -201 1335 -195
rect 1341 -201 1347 -195
rect 1353 -201 1359 -195
rect 1365 -201 1371 -195
rect 1377 -201 1383 -195
rect 1389 -201 1395 -195
rect 1401 -201 1407 -195
rect 1413 -201 1419 -195
rect 1425 -201 1431 -195
rect 1437 -201 1443 -195
rect 1449 -201 1455 -195
rect 1461 -201 1563 -195
rect 1569 -201 1575 -195
rect 1581 -201 1587 -195
rect 1593 -201 1599 -195
rect 1605 -201 1611 -195
rect 1617 -201 1623 -195
rect 1629 -201 1632 -195
rect -108 -204 1632 -201
<< via1 >>
rect -33 567 -27 573
rect 15 567 21 573
rect 63 567 69 573
rect 111 567 117 573
rect 159 567 165 573
rect 207 567 213 573
rect 255 567 261 573
rect 303 567 309 573
rect 351 567 357 573
rect 399 567 405 573
rect 447 567 453 573
rect 495 567 501 573
rect 543 567 549 573
rect 591 567 597 573
rect 639 567 645 573
rect 687 567 693 573
rect 735 567 741 573
rect 783 567 789 573
rect 831 567 837 573
rect 879 567 885 573
rect 927 567 933 573
rect 975 567 981 573
rect 1023 567 1029 573
rect 1071 567 1077 573
rect 1119 567 1125 573
rect 1167 567 1173 573
rect 1215 567 1221 573
rect 1263 567 1269 573
rect 1311 567 1317 573
rect 1359 567 1365 573
rect 1407 567 1413 573
rect 1455 567 1461 573
rect 1503 567 1509 573
rect 1551 567 1557 573
rect -57 543 -51 549
rect -57 531 -51 537
rect -57 519 -51 525
rect -9 543 -3 549
rect -9 531 -3 537
rect -9 519 -3 525
rect 15 543 21 549
rect 15 531 21 537
rect 15 519 21 525
rect 39 543 45 549
rect 39 531 45 537
rect 39 519 45 525
rect 63 543 69 549
rect 63 531 69 537
rect 63 519 69 525
rect 87 543 93 549
rect 87 531 93 537
rect 87 519 93 525
rect 111 543 117 549
rect 111 531 117 537
rect 111 519 117 525
rect 135 543 141 549
rect 135 531 141 537
rect 135 519 141 525
rect 159 543 165 549
rect 159 531 165 537
rect 159 519 165 525
rect 183 543 189 549
rect 183 531 189 537
rect 183 519 189 525
rect 207 543 213 549
rect 207 531 213 537
rect 207 519 213 525
rect 231 543 237 549
rect 231 531 237 537
rect 231 519 237 525
rect 255 543 261 549
rect 255 531 261 537
rect 255 519 261 525
rect 279 543 285 549
rect 279 531 285 537
rect 279 519 285 525
rect 303 543 309 549
rect 303 531 309 537
rect 303 519 309 525
rect 327 543 333 549
rect 327 531 333 537
rect 327 519 333 525
rect 351 543 357 549
rect 351 531 357 537
rect 351 519 357 525
rect 375 543 381 549
rect 375 531 381 537
rect 375 519 381 525
rect 399 543 405 549
rect 399 531 405 537
rect 399 519 405 525
rect 423 543 429 549
rect 423 531 429 537
rect 423 519 429 525
rect 447 543 453 549
rect 447 531 453 537
rect 447 519 453 525
rect 471 543 477 549
rect 471 531 477 537
rect 471 519 477 525
rect 495 543 501 549
rect 495 531 501 537
rect 495 519 501 525
rect 519 543 525 549
rect 519 531 525 537
rect 519 519 525 525
rect 543 543 549 549
rect 543 531 549 537
rect 543 519 549 525
rect 567 543 573 549
rect 567 531 573 537
rect 567 519 573 525
rect 591 543 597 549
rect 591 531 597 537
rect 591 519 597 525
rect 615 543 621 549
rect 615 531 621 537
rect 615 519 621 525
rect 639 543 645 549
rect 639 531 645 537
rect 639 519 645 525
rect 663 543 669 549
rect 663 531 669 537
rect 663 519 669 525
rect 687 543 693 549
rect 687 531 693 537
rect 687 519 693 525
rect 711 543 717 549
rect 711 531 717 537
rect 711 519 717 525
rect 735 543 741 549
rect 735 531 741 537
rect 735 519 741 525
rect 759 543 765 549
rect 759 531 765 537
rect 759 519 765 525
rect 783 543 789 549
rect 783 531 789 537
rect 783 519 789 525
rect 807 543 813 549
rect 807 531 813 537
rect 807 519 813 525
rect 831 543 837 549
rect 831 531 837 537
rect 831 519 837 525
rect 855 543 861 549
rect 855 531 861 537
rect 855 519 861 525
rect 879 543 885 549
rect 879 531 885 537
rect 879 519 885 525
rect 903 543 909 549
rect 903 531 909 537
rect 903 519 909 525
rect 927 543 933 549
rect 927 531 933 537
rect 927 519 933 525
rect 951 543 957 549
rect 951 531 957 537
rect 951 519 957 525
rect 975 543 981 549
rect 975 531 981 537
rect 975 519 981 525
rect 999 543 1005 549
rect 999 531 1005 537
rect 999 519 1005 525
rect 1023 543 1029 549
rect 1023 531 1029 537
rect 1023 519 1029 525
rect 1047 543 1053 549
rect 1047 531 1053 537
rect 1047 519 1053 525
rect 1071 543 1077 549
rect 1071 531 1077 537
rect 1071 519 1077 525
rect 1095 543 1101 549
rect 1095 531 1101 537
rect 1095 519 1101 525
rect 1119 543 1125 549
rect 1119 531 1125 537
rect 1119 519 1125 525
rect 1143 543 1149 549
rect 1143 531 1149 537
rect 1143 519 1149 525
rect 1167 543 1173 549
rect 1167 531 1173 537
rect 1167 519 1173 525
rect 1191 543 1197 549
rect 1191 531 1197 537
rect 1191 519 1197 525
rect 1215 543 1221 549
rect 1215 531 1221 537
rect 1215 519 1221 525
rect 1239 543 1245 549
rect 1239 531 1245 537
rect 1239 519 1245 525
rect 1263 543 1269 549
rect 1263 531 1269 537
rect 1263 519 1269 525
rect 1287 543 1293 549
rect 1287 531 1293 537
rect 1287 519 1293 525
rect 1311 543 1317 549
rect 1311 531 1317 537
rect 1311 519 1317 525
rect 1335 543 1341 549
rect 1335 531 1341 537
rect 1335 519 1341 525
rect 1359 543 1365 549
rect 1359 531 1365 537
rect 1359 519 1365 525
rect 1383 543 1389 549
rect 1383 531 1389 537
rect 1383 519 1389 525
rect 1407 543 1413 549
rect 1407 531 1413 537
rect 1407 519 1413 525
rect 1431 543 1437 549
rect 1431 531 1437 537
rect 1431 519 1437 525
rect 1455 543 1461 549
rect 1455 531 1461 537
rect 1455 519 1461 525
rect 1479 543 1485 549
rect 1479 531 1485 537
rect 1479 519 1485 525
rect 1503 543 1509 549
rect 1503 531 1509 537
rect 1503 519 1509 525
rect 1527 543 1533 549
rect 1527 531 1533 537
rect 1527 519 1533 525
rect 1575 543 1581 549
rect 1575 531 1581 537
rect 1575 519 1581 525
rect -81 447 -75 453
rect -33 447 -27 453
rect 15 447 21 453
rect 63 447 69 453
rect 111 447 117 453
rect 159 447 165 453
rect 207 447 213 453
rect 255 447 261 453
rect 303 447 309 453
rect 351 447 357 453
rect 399 447 405 453
rect 447 447 453 453
rect 495 447 501 453
rect 543 447 549 453
rect 591 447 597 453
rect 639 447 645 453
rect 687 447 693 453
rect 735 447 741 453
rect 783 447 789 453
rect 831 447 837 453
rect 879 447 885 453
rect 927 447 933 453
rect 975 447 981 453
rect 1023 447 1029 453
rect 1071 447 1077 453
rect 1119 447 1125 453
rect 1167 447 1173 453
rect 1215 447 1221 453
rect 1263 447 1269 453
rect 1311 447 1317 453
rect 1359 447 1365 453
rect 1407 447 1413 453
rect 1455 447 1461 453
rect 1503 447 1509 453
rect 1551 447 1557 453
rect 1599 447 1605 453
rect -57 423 -51 429
rect -9 423 -3 429
rect -57 411 -51 417
rect -57 399 -51 405
rect 39 423 45 429
rect -9 411 -3 417
rect -9 399 -3 405
rect 15 399 21 405
rect 87 423 93 429
rect 63 399 69 405
rect 135 423 141 429
rect 87 411 93 417
rect 87 399 93 405
rect 111 399 117 405
rect 183 423 189 429
rect 159 399 165 405
rect 183 411 189 417
rect 183 399 189 405
rect 231 399 237 405
rect 279 423 285 429
rect 327 399 333 405
rect 375 423 381 429
rect 375 411 381 417
rect 375 399 381 405
rect 423 399 429 405
rect 471 423 477 429
rect 519 399 525 405
rect 567 423 573 429
rect 615 423 621 429
rect 567 411 573 417
rect 567 399 573 405
rect 591 399 597 405
rect 663 423 669 429
rect 639 399 645 405
rect 711 423 717 429
rect 663 411 669 417
rect 663 399 669 405
rect 687 399 693 405
rect 759 423 765 429
rect 735 399 741 405
rect 807 423 813 429
rect 759 411 765 417
rect 759 399 765 405
rect 783 399 789 405
rect 855 423 861 429
rect 831 399 837 405
rect 903 423 909 429
rect 855 411 861 417
rect 855 399 861 405
rect 879 399 885 405
rect 951 423 957 429
rect 927 399 933 405
rect 951 411 957 417
rect 951 399 957 405
rect 999 399 1005 405
rect 1047 423 1053 429
rect 1095 399 1101 405
rect 1143 423 1149 429
rect 1143 411 1149 417
rect 1143 399 1149 405
rect 1191 399 1197 405
rect 1239 423 1245 429
rect 1287 399 1293 405
rect 1335 423 1341 429
rect 1383 423 1389 429
rect 1335 411 1341 417
rect 1335 399 1341 405
rect 1359 399 1365 405
rect 1431 423 1437 429
rect 1407 399 1413 405
rect 1479 423 1485 429
rect 1431 411 1437 417
rect 1431 399 1437 405
rect 1455 399 1461 405
rect 1527 423 1533 429
rect 1503 399 1509 405
rect 1575 423 1581 429
rect 1527 411 1533 417
rect 1527 399 1533 405
rect 1575 411 1581 417
rect 1575 399 1581 405
rect 15 375 21 381
rect 63 375 69 381
rect 111 375 117 381
rect 159 375 165 381
rect 207 375 213 381
rect 255 375 261 381
rect 303 375 309 381
rect 351 375 357 381
rect 399 375 405 381
rect 447 375 453 381
rect 495 375 501 381
rect 543 375 549 381
rect 591 375 597 381
rect 639 375 645 381
rect 687 375 693 381
rect 735 375 741 381
rect 783 375 789 381
rect 831 375 837 381
rect 879 375 885 381
rect 927 375 933 381
rect 975 375 981 381
rect 1023 375 1029 381
rect 1071 375 1077 381
rect 1119 375 1125 381
rect 1167 375 1173 381
rect 1215 375 1221 381
rect 1263 375 1269 381
rect 1311 375 1317 381
rect 1359 375 1365 381
rect 1407 375 1413 381
rect 1455 375 1461 381
rect 1503 375 1509 381
rect -57 327 -51 333
rect -9 327 -3 333
rect 183 327 189 333
rect 375 327 381 333
rect 567 327 573 333
rect 759 327 765 333
rect 951 327 957 333
rect 1143 327 1149 333
rect 1335 327 1341 333
rect 1527 327 1533 333
rect 1575 327 1581 333
rect -57 87 -51 93
rect -9 87 -3 93
rect 183 87 189 93
rect 375 87 381 93
rect 567 87 573 93
rect 759 87 765 93
rect 951 87 957 93
rect 1143 87 1149 93
rect 1335 87 1341 93
rect 1527 87 1533 93
rect 1575 87 1581 93
rect 15 63 21 69
rect 63 63 69 69
rect 111 63 117 69
rect 159 63 165 69
rect 207 63 213 69
rect 255 63 261 69
rect 303 63 309 69
rect 351 63 357 69
rect 399 63 405 69
rect 447 63 453 69
rect 495 63 501 69
rect 543 63 549 69
rect 591 63 597 69
rect 639 63 645 69
rect 687 63 693 69
rect 735 63 741 69
rect 783 63 789 69
rect 831 63 837 69
rect 879 63 885 69
rect 927 63 933 69
rect 975 63 981 69
rect 1023 63 1029 69
rect 1071 63 1077 69
rect 1119 63 1125 69
rect 1167 63 1173 69
rect 1215 63 1221 69
rect 1263 63 1269 69
rect 1311 63 1317 69
rect 1359 63 1365 69
rect 1407 63 1413 69
rect 1455 63 1461 69
rect 1503 63 1509 69
rect -57 39 -51 45
rect -57 27 -51 33
rect -57 15 -51 21
rect -9 39 -3 45
rect -9 27 -3 33
rect -9 15 -3 21
rect 39 39 45 45
rect 39 27 45 33
rect 39 15 45 21
rect 87 39 93 45
rect 87 27 93 33
rect 87 15 93 21
rect 135 39 141 45
rect 135 27 141 33
rect 135 15 141 21
rect 183 39 189 45
rect 183 27 189 33
rect 183 15 189 21
rect 279 39 285 45
rect 279 27 285 33
rect 279 15 285 21
rect 375 39 381 45
rect 375 27 381 33
rect 375 15 381 21
rect 471 39 477 45
rect 471 27 477 33
rect 471 15 477 21
rect 567 39 573 45
rect 567 27 573 33
rect 567 15 573 21
rect 615 39 621 45
rect 615 27 621 33
rect 615 15 621 21
rect 663 39 669 45
rect 663 27 669 33
rect 663 15 669 21
rect 711 39 717 45
rect 711 27 717 33
rect 711 15 717 21
rect 759 39 765 45
rect 759 27 765 33
rect 759 15 765 21
rect 807 39 813 45
rect 807 27 813 33
rect 807 15 813 21
rect 855 39 861 45
rect 855 27 861 33
rect 855 15 861 21
rect 903 39 909 45
rect 903 27 909 33
rect 903 15 909 21
rect 951 39 957 45
rect 951 27 957 33
rect 951 15 957 21
rect 1047 39 1053 45
rect 1047 27 1053 33
rect 1047 15 1053 21
rect 1143 39 1149 45
rect 1143 27 1149 33
rect 1143 15 1149 21
rect 1239 39 1245 45
rect 1239 27 1245 33
rect 1239 15 1245 21
rect 1335 39 1341 45
rect 1335 27 1341 33
rect 1335 15 1341 21
rect 1383 39 1389 45
rect 1383 27 1389 33
rect 1383 15 1389 21
rect 1431 39 1437 45
rect 1431 27 1437 33
rect 1431 15 1437 21
rect 1479 39 1485 45
rect 1479 27 1485 33
rect 1479 15 1485 21
rect 1527 39 1533 45
rect 1527 27 1533 33
rect 1527 15 1533 21
rect 1575 39 1581 45
rect 1575 27 1581 33
rect 1575 15 1581 21
rect -57 -9 -51 -3
rect -9 -9 -3 -3
rect 183 -9 189 -3
rect 375 -9 381 -3
rect 567 -9 573 -3
rect 759 -9 765 -3
rect 951 -9 957 -3
rect 1143 -9 1149 -3
rect 1335 -9 1341 -3
rect 1527 -9 1533 -3
rect 1575 -9 1581 -3
<< metal2 >>
rect -84 597 -72 600
rect -84 591 -81 597
rect -75 591 -72 597
rect -84 549 -72 591
rect 1596 597 1608 600
rect 1596 591 1599 597
rect 1605 591 1608 597
rect -36 573 -24 576
rect -36 567 -33 573
rect -27 567 -24 573
rect -36 564 -24 567
rect 12 573 24 576
rect 12 567 15 573
rect 21 567 24 573
rect 12 564 24 567
rect 60 573 72 576
rect 60 567 63 573
rect 69 567 72 573
rect 60 564 72 567
rect 108 573 120 576
rect 108 567 111 573
rect 117 567 120 573
rect 108 564 120 567
rect 156 573 168 576
rect 156 567 159 573
rect 165 567 168 573
rect 156 564 168 567
rect 204 573 216 576
rect 204 567 207 573
rect 213 567 216 573
rect 204 564 216 567
rect 252 573 264 576
rect 252 567 255 573
rect 261 567 264 573
rect 252 564 264 567
rect 300 573 312 576
rect 300 567 303 573
rect 309 567 312 573
rect 300 564 312 567
rect 348 573 360 576
rect 348 567 351 573
rect 357 567 360 573
rect 348 564 360 567
rect 396 573 408 576
rect 396 567 399 573
rect 405 567 408 573
rect 396 564 408 567
rect 444 573 456 576
rect 444 567 447 573
rect 453 567 456 573
rect 444 564 456 567
rect 492 573 504 576
rect 492 567 495 573
rect 501 567 504 573
rect 492 564 504 567
rect 540 573 552 576
rect 540 567 543 573
rect 549 567 552 573
rect 540 564 552 567
rect 588 573 600 576
rect 588 567 591 573
rect 597 567 600 573
rect 588 564 600 567
rect 636 573 648 576
rect 636 567 639 573
rect 645 567 648 573
rect 636 564 648 567
rect 684 573 696 576
rect 684 567 687 573
rect 693 567 696 573
rect 684 564 696 567
rect 732 573 744 576
rect 732 567 735 573
rect 741 567 744 573
rect 732 564 744 567
rect 780 573 792 576
rect 780 567 783 573
rect 789 567 792 573
rect 780 564 792 567
rect 828 573 840 576
rect 828 567 831 573
rect 837 567 840 573
rect 828 564 840 567
rect 876 573 888 576
rect 876 567 879 573
rect 885 567 888 573
rect 876 564 888 567
rect 924 573 936 576
rect 924 567 927 573
rect 933 567 936 573
rect 924 564 936 567
rect 972 573 984 576
rect 972 567 975 573
rect 981 567 984 573
rect 972 564 984 567
rect 1020 573 1032 576
rect 1020 567 1023 573
rect 1029 567 1032 573
rect 1020 564 1032 567
rect 1068 573 1080 576
rect 1068 567 1071 573
rect 1077 567 1080 573
rect 1068 564 1080 567
rect 1116 573 1128 576
rect 1116 567 1119 573
rect 1125 567 1128 573
rect 1116 564 1128 567
rect 1164 573 1176 576
rect 1164 567 1167 573
rect 1173 567 1176 573
rect 1164 564 1176 567
rect 1212 573 1224 576
rect 1212 567 1215 573
rect 1221 567 1224 573
rect 1212 564 1224 567
rect 1260 573 1272 576
rect 1260 567 1263 573
rect 1269 567 1272 573
rect 1260 564 1272 567
rect 1308 573 1320 576
rect 1308 567 1311 573
rect 1317 567 1320 573
rect 1308 564 1320 567
rect 1356 573 1368 576
rect 1356 567 1359 573
rect 1365 567 1368 573
rect 1356 564 1368 567
rect 1404 573 1416 576
rect 1404 567 1407 573
rect 1413 567 1416 573
rect 1404 564 1416 567
rect 1452 573 1464 576
rect 1452 567 1455 573
rect 1461 567 1464 573
rect 1452 564 1464 567
rect 1500 573 1512 576
rect 1500 567 1503 573
rect 1509 567 1512 573
rect 1500 564 1512 567
rect 1548 573 1560 576
rect 1548 567 1551 573
rect 1557 567 1560 573
rect 1548 564 1560 567
rect -84 543 -81 549
rect -75 543 -72 549
rect -84 537 -72 543
rect -84 531 -81 537
rect -75 531 -72 537
rect -84 525 -72 531
rect -84 519 -81 525
rect -75 519 -72 525
rect -84 516 -72 519
rect -60 549 -48 552
rect -60 543 -57 549
rect -51 543 -48 549
rect -60 537 -48 543
rect -60 531 -57 537
rect -51 531 -48 537
rect -60 525 -48 531
rect -60 519 -57 525
rect -51 519 -48 525
rect -60 477 -48 519
rect -60 471 -57 477
rect -51 471 -48 477
rect -84 453 -72 456
rect -84 447 -81 453
rect -75 447 -72 453
rect -84 444 -72 447
rect -60 429 -48 471
rect -12 549 0 552
rect -12 543 -9 549
rect -3 543 0 549
rect -12 537 0 543
rect -12 531 -9 537
rect -3 531 0 537
rect -12 525 0 531
rect -12 519 -9 525
rect -3 519 0 525
rect -12 477 0 519
rect 12 549 24 552
rect 12 543 15 549
rect 21 543 24 549
rect 12 537 24 543
rect 12 531 15 537
rect 21 531 24 537
rect 12 525 24 531
rect 12 519 15 525
rect 21 519 24 525
rect 12 516 24 519
rect 36 549 48 552
rect 36 543 39 549
rect 45 543 48 549
rect 36 537 48 543
rect 36 531 39 537
rect 45 531 48 537
rect 36 525 48 531
rect 36 519 39 525
rect 45 519 48 525
rect -12 471 -9 477
rect -3 471 0 477
rect -36 453 -24 456
rect -36 447 -33 453
rect -27 447 -24 453
rect -36 444 -24 447
rect -60 423 -57 429
rect -51 423 -48 429
rect -60 417 -48 423
rect -60 411 -57 417
rect -51 411 -48 417
rect -60 405 -48 411
rect -60 399 -57 405
rect -51 399 -48 405
rect -60 396 -48 399
rect -12 432 0 471
rect 36 477 48 519
rect 60 549 72 552
rect 60 543 63 549
rect 69 543 72 549
rect 60 537 72 543
rect 60 531 63 537
rect 69 531 72 537
rect 60 525 72 531
rect 60 519 63 525
rect 69 519 72 525
rect 60 516 72 519
rect 84 549 96 552
rect 84 543 87 549
rect 93 543 96 549
rect 84 537 96 543
rect 84 531 87 537
rect 93 531 96 537
rect 84 525 96 531
rect 84 519 87 525
rect 93 519 96 525
rect 36 471 39 477
rect 45 471 48 477
rect 12 453 24 456
rect 12 447 15 453
rect 21 447 24 453
rect 12 444 24 447
rect 36 432 48 471
rect 84 477 96 519
rect 108 549 120 552
rect 108 543 111 549
rect 117 543 120 549
rect 108 537 120 543
rect 108 531 111 537
rect 117 531 120 537
rect 108 525 120 531
rect 108 519 111 525
rect 117 519 120 525
rect 108 516 120 519
rect 132 549 144 552
rect 132 543 135 549
rect 141 543 144 549
rect 132 537 144 543
rect 132 531 135 537
rect 141 531 144 537
rect 132 525 144 531
rect 132 519 135 525
rect 141 519 144 525
rect 84 471 87 477
rect 93 471 96 477
rect 60 453 72 456
rect 60 447 63 453
rect 69 447 72 453
rect 60 444 72 447
rect 84 432 96 471
rect 132 477 144 519
rect 156 549 168 552
rect 156 543 159 549
rect 165 543 168 549
rect 156 537 168 543
rect 156 531 159 537
rect 165 531 168 537
rect 156 525 168 531
rect 156 519 159 525
rect 165 519 168 525
rect 156 516 168 519
rect 180 549 192 552
rect 180 543 183 549
rect 189 543 192 549
rect 180 537 192 543
rect 180 531 183 537
rect 189 531 192 537
rect 180 525 192 531
rect 180 519 183 525
rect 189 519 192 525
rect 132 471 135 477
rect 141 471 144 477
rect 108 453 120 456
rect 108 447 111 453
rect 117 447 120 453
rect 108 444 120 447
rect 132 432 144 471
rect 180 477 192 519
rect 204 549 216 552
rect 204 543 207 549
rect 213 543 216 549
rect 204 537 216 543
rect 204 531 207 537
rect 213 531 216 537
rect 204 525 216 531
rect 204 519 207 525
rect 213 519 216 525
rect 204 516 216 519
rect 228 549 240 552
rect 228 543 231 549
rect 237 543 240 549
rect 228 537 240 543
rect 228 531 231 537
rect 237 531 240 537
rect 228 525 240 531
rect 228 519 231 525
rect 237 519 240 525
rect 180 471 183 477
rect 189 471 192 477
rect 156 453 168 456
rect 156 447 159 453
rect 165 447 168 453
rect 156 444 168 447
rect 180 432 192 471
rect 228 477 240 519
rect 252 549 264 552
rect 252 543 255 549
rect 261 543 264 549
rect 252 537 264 543
rect 252 531 255 537
rect 261 531 264 537
rect 252 525 264 531
rect 252 519 255 525
rect 261 519 264 525
rect 252 516 264 519
rect 276 549 288 552
rect 276 543 279 549
rect 285 543 288 549
rect 276 537 288 543
rect 276 531 279 537
rect 285 531 288 537
rect 276 525 288 531
rect 276 519 279 525
rect 285 519 288 525
rect 228 471 231 477
rect 237 471 240 477
rect 204 453 216 456
rect 204 447 207 453
rect 213 447 216 453
rect 204 444 216 447
rect 228 432 240 471
rect 276 477 288 519
rect 300 549 312 552
rect 300 543 303 549
rect 309 543 312 549
rect 300 537 312 543
rect 300 531 303 537
rect 309 531 312 537
rect 300 525 312 531
rect 300 519 303 525
rect 309 519 312 525
rect 300 516 312 519
rect 324 549 336 552
rect 324 543 327 549
rect 333 543 336 549
rect 324 537 336 543
rect 324 531 327 537
rect 333 531 336 537
rect 324 525 336 531
rect 324 519 327 525
rect 333 519 336 525
rect 276 471 279 477
rect 285 471 288 477
rect 252 453 264 456
rect 252 447 255 453
rect 261 447 264 453
rect 252 444 264 447
rect 276 432 288 471
rect 324 477 336 519
rect 348 549 360 552
rect 348 543 351 549
rect 357 543 360 549
rect 348 537 360 543
rect 348 531 351 537
rect 357 531 360 537
rect 348 525 360 531
rect 348 519 351 525
rect 357 519 360 525
rect 348 516 360 519
rect 372 549 384 552
rect 372 543 375 549
rect 381 543 384 549
rect 372 537 384 543
rect 372 531 375 537
rect 381 531 384 537
rect 372 525 384 531
rect 372 519 375 525
rect 381 519 384 525
rect 324 471 327 477
rect 333 471 336 477
rect 300 453 312 456
rect 300 447 303 453
rect 309 447 312 453
rect 300 444 312 447
rect 324 444 336 471
rect 372 477 384 519
rect 396 549 408 552
rect 396 543 399 549
rect 405 543 408 549
rect 396 537 408 543
rect 396 531 399 537
rect 405 531 408 537
rect 396 525 408 531
rect 396 519 399 525
rect 405 519 408 525
rect 396 516 408 519
rect 420 549 432 552
rect 420 543 423 549
rect 429 543 432 549
rect 420 537 432 543
rect 420 531 423 537
rect 429 531 432 537
rect 420 525 432 531
rect 420 519 423 525
rect 429 519 432 525
rect 372 471 375 477
rect 381 471 384 477
rect 348 453 360 456
rect 348 447 351 453
rect 357 447 360 453
rect 348 444 360 447
rect 372 432 384 471
rect 420 477 432 519
rect 444 549 456 552
rect 444 543 447 549
rect 453 543 456 549
rect 444 537 456 543
rect 444 531 447 537
rect 453 531 456 537
rect 444 525 456 531
rect 444 519 447 525
rect 453 519 456 525
rect 444 516 456 519
rect 468 549 480 552
rect 468 543 471 549
rect 477 543 480 549
rect 468 537 480 543
rect 468 531 471 537
rect 477 531 480 537
rect 468 525 480 531
rect 468 519 471 525
rect 477 519 480 525
rect 420 471 423 477
rect 429 471 432 477
rect 396 453 408 456
rect 396 447 399 453
rect 405 447 408 453
rect 396 444 408 447
rect 420 432 432 471
rect 468 477 480 519
rect 492 549 504 552
rect 492 543 495 549
rect 501 543 504 549
rect 492 537 504 543
rect 492 531 495 537
rect 501 531 504 537
rect 492 525 504 531
rect 492 519 495 525
rect 501 519 504 525
rect 492 516 504 519
rect 516 549 528 552
rect 516 543 519 549
rect 525 543 528 549
rect 516 537 528 543
rect 516 531 519 537
rect 525 531 528 537
rect 516 525 528 531
rect 516 519 519 525
rect 525 519 528 525
rect 468 471 471 477
rect 477 471 480 477
rect 444 453 456 456
rect 444 447 447 453
rect 453 447 456 453
rect 444 444 456 447
rect 468 432 480 471
rect 516 477 528 519
rect 540 549 552 552
rect 540 543 543 549
rect 549 543 552 549
rect 540 537 552 543
rect 540 531 543 537
rect 549 531 552 537
rect 540 525 552 531
rect 540 519 543 525
rect 549 519 552 525
rect 540 516 552 519
rect 564 549 576 552
rect 564 543 567 549
rect 573 543 576 549
rect 564 537 576 543
rect 564 531 567 537
rect 573 531 576 537
rect 564 525 576 531
rect 564 519 567 525
rect 573 519 576 525
rect 516 471 519 477
rect 525 471 528 477
rect 492 453 504 456
rect 492 447 495 453
rect 501 447 504 453
rect 492 444 504 447
rect 516 444 528 471
rect 564 477 576 519
rect 588 549 600 552
rect 588 543 591 549
rect 597 543 600 549
rect 588 537 600 543
rect 588 531 591 537
rect 597 531 600 537
rect 588 525 600 531
rect 588 519 591 525
rect 597 519 600 525
rect 588 516 600 519
rect 612 549 624 552
rect 612 543 615 549
rect 621 543 624 549
rect 612 537 624 543
rect 612 531 615 537
rect 621 531 624 537
rect 612 525 624 531
rect 612 519 615 525
rect 621 519 624 525
rect 564 471 567 477
rect 573 471 576 477
rect 540 453 552 456
rect 540 447 543 453
rect 549 447 552 453
rect 540 444 552 447
rect 564 432 576 471
rect 612 477 624 519
rect 636 549 648 552
rect 636 543 639 549
rect 645 543 648 549
rect 636 537 648 543
rect 636 531 639 537
rect 645 531 648 537
rect 636 525 648 531
rect 636 519 639 525
rect 645 519 648 525
rect 636 516 648 519
rect 660 549 672 552
rect 660 543 663 549
rect 669 543 672 549
rect 660 537 672 543
rect 660 531 663 537
rect 669 531 672 537
rect 660 525 672 531
rect 660 519 663 525
rect 669 519 672 525
rect 612 471 615 477
rect 621 471 624 477
rect 588 453 600 456
rect 588 447 591 453
rect 597 447 600 453
rect 588 444 600 447
rect 612 432 624 471
rect 660 477 672 519
rect 684 549 696 552
rect 684 543 687 549
rect 693 543 696 549
rect 684 537 696 543
rect 684 531 687 537
rect 693 531 696 537
rect 684 525 696 531
rect 684 519 687 525
rect 693 519 696 525
rect 684 516 696 519
rect 708 549 720 552
rect 708 543 711 549
rect 717 543 720 549
rect 708 537 720 543
rect 708 531 711 537
rect 717 531 720 537
rect 708 525 720 531
rect 708 519 711 525
rect 717 519 720 525
rect 660 471 663 477
rect 669 471 672 477
rect 636 453 648 456
rect 636 447 639 453
rect 645 447 648 453
rect 636 444 648 447
rect 660 432 672 471
rect 708 477 720 519
rect 732 549 744 552
rect 732 543 735 549
rect 741 543 744 549
rect 732 537 744 543
rect 732 531 735 537
rect 741 531 744 537
rect 732 525 744 531
rect 732 519 735 525
rect 741 519 744 525
rect 732 516 744 519
rect 756 549 768 552
rect 756 543 759 549
rect 765 543 768 549
rect 756 537 768 543
rect 756 531 759 537
rect 765 531 768 537
rect 756 525 768 531
rect 756 519 759 525
rect 765 519 768 525
rect 708 471 711 477
rect 717 471 720 477
rect 684 453 696 456
rect 684 447 687 453
rect 693 447 696 453
rect 684 444 696 447
rect 708 432 720 471
rect 756 477 768 519
rect 780 549 792 552
rect 780 543 783 549
rect 789 543 792 549
rect 780 537 792 543
rect 780 531 783 537
rect 789 531 792 537
rect 780 525 792 531
rect 780 519 783 525
rect 789 519 792 525
rect 780 516 792 519
rect 804 549 816 552
rect 804 543 807 549
rect 813 543 816 549
rect 804 537 816 543
rect 804 531 807 537
rect 813 531 816 537
rect 804 525 816 531
rect 804 519 807 525
rect 813 519 816 525
rect 756 471 759 477
rect 765 471 768 477
rect 732 453 744 456
rect 732 447 735 453
rect 741 447 744 453
rect 732 444 744 447
rect 756 432 768 471
rect 804 477 816 519
rect 828 549 840 552
rect 828 543 831 549
rect 837 543 840 549
rect 828 537 840 543
rect 828 531 831 537
rect 837 531 840 537
rect 828 525 840 531
rect 828 519 831 525
rect 837 519 840 525
rect 828 516 840 519
rect 852 549 864 552
rect 852 543 855 549
rect 861 543 864 549
rect 852 537 864 543
rect 852 531 855 537
rect 861 531 864 537
rect 852 525 864 531
rect 852 519 855 525
rect 861 519 864 525
rect 804 471 807 477
rect 813 471 816 477
rect 780 453 792 456
rect 780 447 783 453
rect 789 447 792 453
rect 780 444 792 447
rect 804 432 816 471
rect 852 477 864 519
rect 876 549 888 552
rect 876 543 879 549
rect 885 543 888 549
rect 876 537 888 543
rect 876 531 879 537
rect 885 531 888 537
rect 876 525 888 531
rect 876 519 879 525
rect 885 519 888 525
rect 876 516 888 519
rect 900 549 912 552
rect 900 543 903 549
rect 909 543 912 549
rect 900 537 912 543
rect 900 531 903 537
rect 909 531 912 537
rect 900 525 912 531
rect 900 519 903 525
rect 909 519 912 525
rect 852 471 855 477
rect 861 471 864 477
rect 828 453 840 456
rect 828 447 831 453
rect 837 447 840 453
rect 828 444 840 447
rect 852 432 864 471
rect 900 477 912 519
rect 924 549 936 552
rect 924 543 927 549
rect 933 543 936 549
rect 924 537 936 543
rect 924 531 927 537
rect 933 531 936 537
rect 924 525 936 531
rect 924 519 927 525
rect 933 519 936 525
rect 924 516 936 519
rect 948 549 960 552
rect 948 543 951 549
rect 957 543 960 549
rect 948 537 960 543
rect 948 531 951 537
rect 957 531 960 537
rect 948 525 960 531
rect 948 519 951 525
rect 957 519 960 525
rect 900 471 903 477
rect 909 471 912 477
rect 876 453 888 456
rect 876 447 879 453
rect 885 447 888 453
rect 876 444 888 447
rect 900 432 912 471
rect 948 477 960 519
rect 972 549 984 552
rect 972 543 975 549
rect 981 543 984 549
rect 972 537 984 543
rect 972 531 975 537
rect 981 531 984 537
rect 972 525 984 531
rect 972 519 975 525
rect 981 519 984 525
rect 972 516 984 519
rect 996 549 1008 552
rect 996 543 999 549
rect 1005 543 1008 549
rect 996 537 1008 543
rect 996 531 999 537
rect 1005 531 1008 537
rect 996 525 1008 531
rect 996 519 999 525
rect 1005 519 1008 525
rect 948 471 951 477
rect 957 471 960 477
rect 924 453 936 456
rect 924 447 927 453
rect 933 447 936 453
rect 924 444 936 447
rect 948 432 960 471
rect 996 477 1008 519
rect 1020 549 1032 552
rect 1020 543 1023 549
rect 1029 543 1032 549
rect 1020 537 1032 543
rect 1020 531 1023 537
rect 1029 531 1032 537
rect 1020 525 1032 531
rect 1020 519 1023 525
rect 1029 519 1032 525
rect 1020 516 1032 519
rect 1044 549 1056 552
rect 1044 543 1047 549
rect 1053 543 1056 549
rect 1044 537 1056 543
rect 1044 531 1047 537
rect 1053 531 1056 537
rect 1044 525 1056 531
rect 1044 519 1047 525
rect 1053 519 1056 525
rect 996 471 999 477
rect 1005 471 1008 477
rect 972 453 984 456
rect 972 447 975 453
rect 981 447 984 453
rect 972 444 984 447
rect 996 444 1008 471
rect 1044 477 1056 519
rect 1068 549 1080 552
rect 1068 543 1071 549
rect 1077 543 1080 549
rect 1068 537 1080 543
rect 1068 531 1071 537
rect 1077 531 1080 537
rect 1068 525 1080 531
rect 1068 519 1071 525
rect 1077 519 1080 525
rect 1068 516 1080 519
rect 1092 549 1104 552
rect 1092 543 1095 549
rect 1101 543 1104 549
rect 1092 537 1104 543
rect 1092 531 1095 537
rect 1101 531 1104 537
rect 1092 525 1104 531
rect 1092 519 1095 525
rect 1101 519 1104 525
rect 1044 471 1047 477
rect 1053 471 1056 477
rect 1020 453 1032 456
rect 1020 447 1023 453
rect 1029 447 1032 453
rect 1020 444 1032 447
rect 1044 432 1056 471
rect 1092 477 1104 519
rect 1116 549 1128 552
rect 1116 543 1119 549
rect 1125 543 1128 549
rect 1116 537 1128 543
rect 1116 531 1119 537
rect 1125 531 1128 537
rect 1116 525 1128 531
rect 1116 519 1119 525
rect 1125 519 1128 525
rect 1116 516 1128 519
rect 1140 549 1152 552
rect 1140 543 1143 549
rect 1149 543 1152 549
rect 1140 537 1152 543
rect 1140 531 1143 537
rect 1149 531 1152 537
rect 1140 525 1152 531
rect 1140 519 1143 525
rect 1149 519 1152 525
rect 1092 471 1095 477
rect 1101 471 1104 477
rect 1068 453 1080 456
rect 1068 447 1071 453
rect 1077 447 1080 453
rect 1068 444 1080 447
rect 1092 432 1104 471
rect 1140 477 1152 519
rect 1164 549 1176 552
rect 1164 543 1167 549
rect 1173 543 1176 549
rect 1164 537 1176 543
rect 1164 531 1167 537
rect 1173 531 1176 537
rect 1164 525 1176 531
rect 1164 519 1167 525
rect 1173 519 1176 525
rect 1164 516 1176 519
rect 1188 549 1200 552
rect 1188 543 1191 549
rect 1197 543 1200 549
rect 1188 537 1200 543
rect 1188 531 1191 537
rect 1197 531 1200 537
rect 1188 525 1200 531
rect 1188 519 1191 525
rect 1197 519 1200 525
rect 1140 471 1143 477
rect 1149 471 1152 477
rect 1116 453 1128 456
rect 1116 447 1119 453
rect 1125 447 1128 453
rect 1116 444 1128 447
rect 1140 432 1152 471
rect 1188 477 1200 519
rect 1212 549 1224 552
rect 1212 543 1215 549
rect 1221 543 1224 549
rect 1212 537 1224 543
rect 1212 531 1215 537
rect 1221 531 1224 537
rect 1212 525 1224 531
rect 1212 519 1215 525
rect 1221 519 1224 525
rect 1212 516 1224 519
rect 1236 549 1248 552
rect 1236 543 1239 549
rect 1245 543 1248 549
rect 1236 537 1248 543
rect 1236 531 1239 537
rect 1245 531 1248 537
rect 1236 525 1248 531
rect 1236 519 1239 525
rect 1245 519 1248 525
rect 1188 471 1191 477
rect 1197 471 1200 477
rect 1164 453 1176 456
rect 1164 447 1167 453
rect 1173 447 1176 453
rect 1164 444 1176 447
rect 1188 444 1200 471
rect 1236 477 1248 519
rect 1260 549 1272 552
rect 1260 543 1263 549
rect 1269 543 1272 549
rect 1260 537 1272 543
rect 1260 531 1263 537
rect 1269 531 1272 537
rect 1260 525 1272 531
rect 1260 519 1263 525
rect 1269 519 1272 525
rect 1260 516 1272 519
rect 1284 549 1296 552
rect 1284 543 1287 549
rect 1293 543 1296 549
rect 1284 537 1296 543
rect 1284 531 1287 537
rect 1293 531 1296 537
rect 1284 525 1296 531
rect 1284 519 1287 525
rect 1293 519 1296 525
rect 1236 471 1239 477
rect 1245 471 1248 477
rect 1212 453 1224 456
rect 1212 447 1215 453
rect 1221 447 1224 453
rect 1212 444 1224 447
rect 1236 432 1248 471
rect 1284 477 1296 519
rect 1308 549 1320 552
rect 1308 543 1311 549
rect 1317 543 1320 549
rect 1308 537 1320 543
rect 1308 531 1311 537
rect 1317 531 1320 537
rect 1308 525 1320 531
rect 1308 519 1311 525
rect 1317 519 1320 525
rect 1308 516 1320 519
rect 1332 549 1344 552
rect 1332 543 1335 549
rect 1341 543 1344 549
rect 1332 537 1344 543
rect 1332 531 1335 537
rect 1341 531 1344 537
rect 1332 525 1344 531
rect 1332 519 1335 525
rect 1341 519 1344 525
rect 1284 471 1287 477
rect 1293 471 1296 477
rect 1260 453 1272 456
rect 1260 447 1263 453
rect 1269 447 1272 453
rect 1260 444 1272 447
rect 1284 432 1296 471
rect 1332 477 1344 519
rect 1356 549 1368 552
rect 1356 543 1359 549
rect 1365 543 1368 549
rect 1356 537 1368 543
rect 1356 531 1359 537
rect 1365 531 1368 537
rect 1356 525 1368 531
rect 1356 519 1359 525
rect 1365 519 1368 525
rect 1356 516 1368 519
rect 1380 549 1392 552
rect 1380 543 1383 549
rect 1389 543 1392 549
rect 1380 537 1392 543
rect 1380 531 1383 537
rect 1389 531 1392 537
rect 1380 525 1392 531
rect 1380 519 1383 525
rect 1389 519 1392 525
rect 1332 471 1335 477
rect 1341 471 1344 477
rect 1308 453 1320 456
rect 1308 447 1311 453
rect 1317 447 1320 453
rect 1308 444 1320 447
rect 1332 432 1344 471
rect 1380 477 1392 519
rect 1404 549 1416 552
rect 1404 543 1407 549
rect 1413 543 1416 549
rect 1404 537 1416 543
rect 1404 531 1407 537
rect 1413 531 1416 537
rect 1404 525 1416 531
rect 1404 519 1407 525
rect 1413 519 1416 525
rect 1404 516 1416 519
rect 1428 549 1440 552
rect 1428 543 1431 549
rect 1437 543 1440 549
rect 1428 537 1440 543
rect 1428 531 1431 537
rect 1437 531 1440 537
rect 1428 525 1440 531
rect 1428 519 1431 525
rect 1437 519 1440 525
rect 1380 471 1383 477
rect 1389 471 1392 477
rect 1356 453 1368 456
rect 1356 447 1359 453
rect 1365 447 1368 453
rect 1356 444 1368 447
rect 1380 432 1392 471
rect 1428 477 1440 519
rect 1452 549 1464 552
rect 1452 543 1455 549
rect 1461 543 1464 549
rect 1452 537 1464 543
rect 1452 531 1455 537
rect 1461 531 1464 537
rect 1452 525 1464 531
rect 1452 519 1455 525
rect 1461 519 1464 525
rect 1452 516 1464 519
rect 1476 549 1488 552
rect 1476 543 1479 549
rect 1485 543 1488 549
rect 1476 537 1488 543
rect 1476 531 1479 537
rect 1485 531 1488 537
rect 1476 525 1488 531
rect 1476 519 1479 525
rect 1485 519 1488 525
rect 1428 471 1431 477
rect 1437 471 1440 477
rect 1404 453 1416 456
rect 1404 447 1407 453
rect 1413 447 1416 453
rect 1404 444 1416 447
rect 1428 432 1440 471
rect 1476 477 1488 519
rect 1500 549 1512 552
rect 1500 543 1503 549
rect 1509 543 1512 549
rect 1500 537 1512 543
rect 1500 531 1503 537
rect 1509 531 1512 537
rect 1500 525 1512 531
rect 1500 519 1503 525
rect 1509 519 1512 525
rect 1500 516 1512 519
rect 1524 549 1536 552
rect 1524 543 1527 549
rect 1533 543 1536 549
rect 1524 537 1536 543
rect 1524 531 1527 537
rect 1533 531 1536 537
rect 1524 525 1536 531
rect 1524 519 1527 525
rect 1533 519 1536 525
rect 1476 471 1479 477
rect 1485 471 1488 477
rect 1452 453 1464 456
rect 1452 447 1455 453
rect 1461 447 1464 453
rect 1452 444 1464 447
rect 1476 432 1488 471
rect 1524 477 1536 519
rect 1524 471 1527 477
rect 1533 471 1536 477
rect 1500 453 1512 456
rect 1500 447 1503 453
rect 1509 447 1512 453
rect 1500 444 1512 447
rect 1524 432 1536 471
rect 1572 549 1584 552
rect 1572 543 1575 549
rect 1581 543 1584 549
rect 1572 537 1584 543
rect 1572 531 1575 537
rect 1581 531 1584 537
rect 1572 525 1584 531
rect 1572 519 1575 525
rect 1581 519 1584 525
rect 1572 477 1584 519
rect 1596 549 1608 591
rect 1596 543 1599 549
rect 1605 543 1608 549
rect 1596 537 1608 543
rect 1596 531 1599 537
rect 1605 531 1608 537
rect 1596 525 1608 531
rect 1596 519 1599 525
rect 1605 519 1608 525
rect 1596 516 1608 519
rect 1572 471 1575 477
rect 1581 471 1584 477
rect 1548 453 1560 456
rect 1548 447 1551 453
rect 1557 447 1560 453
rect 1548 444 1560 447
rect -12 429 1536 432
rect -12 423 -9 429
rect -3 423 39 429
rect 45 423 87 429
rect 93 423 135 429
rect 141 423 183 429
rect 189 423 279 429
rect 285 423 375 429
rect 381 423 471 429
rect 477 423 567 429
rect 573 423 615 429
rect 621 423 663 429
rect 669 423 711 429
rect 717 423 759 429
rect 765 423 807 429
rect 813 423 855 429
rect 861 423 903 429
rect 909 423 951 429
rect 957 423 1047 429
rect 1053 423 1143 429
rect 1149 423 1239 429
rect 1245 423 1335 429
rect 1341 423 1383 429
rect 1389 423 1431 429
rect 1437 423 1479 429
rect 1485 423 1527 429
rect 1533 423 1536 429
rect -12 420 1536 423
rect -12 417 0 420
rect -12 411 -9 417
rect -3 411 0 417
rect -12 405 0 411
rect 84 417 96 420
rect 84 411 87 417
rect 93 411 96 417
rect -12 399 -9 405
rect -3 399 0 405
rect -12 396 0 399
rect 12 405 72 408
rect 12 399 15 405
rect 21 399 63 405
rect 69 399 72 405
rect 12 396 72 399
rect 84 405 96 411
rect 180 417 192 420
rect 180 411 183 417
rect 189 411 192 417
rect 84 399 87 405
rect 93 399 96 405
rect 84 396 96 399
rect 108 405 168 408
rect 108 399 111 405
rect 117 399 159 405
rect 165 399 168 405
rect 108 396 168 399
rect 180 405 192 411
rect 372 417 384 420
rect 372 411 375 417
rect 381 411 384 417
rect 180 399 183 405
rect 189 399 192 405
rect 180 396 192 399
rect 228 405 336 408
rect 228 399 231 405
rect 237 399 327 405
rect 333 399 336 405
rect 228 396 336 399
rect 372 405 384 411
rect 564 417 576 420
rect 564 411 567 417
rect 573 411 576 417
rect 372 399 375 405
rect 381 399 384 405
rect 372 396 384 399
rect 420 405 528 408
rect 420 399 423 405
rect 429 399 519 405
rect 525 399 528 405
rect 420 396 528 399
rect 564 405 576 411
rect 660 417 672 420
rect 660 411 663 417
rect 669 411 672 417
rect 564 399 567 405
rect 573 399 576 405
rect 564 396 576 399
rect 588 405 648 408
rect 588 399 591 405
rect 597 399 639 405
rect 645 399 648 405
rect 588 396 648 399
rect 660 405 672 411
rect 756 417 768 420
rect 756 411 759 417
rect 765 411 768 417
rect 660 399 663 405
rect 669 399 672 405
rect 660 396 672 399
rect 684 405 744 408
rect 684 399 687 405
rect 693 399 735 405
rect 741 399 744 405
rect 684 396 744 399
rect 756 405 768 411
rect 852 417 864 420
rect 852 411 855 417
rect 861 411 864 417
rect 756 399 759 405
rect 765 399 768 405
rect 756 396 768 399
rect 780 405 840 408
rect 780 399 783 405
rect 789 399 831 405
rect 837 399 840 405
rect 780 396 840 399
rect 852 405 864 411
rect 948 417 960 420
rect 948 411 951 417
rect 957 411 960 417
rect 852 399 855 405
rect 861 399 864 405
rect 852 396 864 399
rect 876 405 936 408
rect 876 399 879 405
rect 885 399 927 405
rect 933 399 936 405
rect 876 396 936 399
rect 948 405 960 411
rect 1140 417 1152 420
rect 1140 411 1143 417
rect 1149 411 1152 417
rect 948 399 951 405
rect 957 399 960 405
rect 948 396 960 399
rect 996 405 1104 408
rect 996 399 999 405
rect 1005 399 1095 405
rect 1101 399 1104 405
rect 996 396 1104 399
rect 1140 405 1152 411
rect 1332 417 1344 420
rect 1332 411 1335 417
rect 1341 411 1344 417
rect 1140 399 1143 405
rect 1149 399 1152 405
rect 1140 396 1152 399
rect 1188 405 1296 408
rect 1188 399 1191 405
rect 1197 399 1287 405
rect 1293 399 1296 405
rect 1188 396 1296 399
rect 1332 405 1344 411
rect 1428 417 1440 420
rect 1428 411 1431 417
rect 1437 411 1440 417
rect 1332 399 1335 405
rect 1341 399 1344 405
rect 1332 396 1344 399
rect 1356 405 1416 408
rect 1356 399 1359 405
rect 1365 399 1407 405
rect 1413 399 1416 405
rect 1356 396 1416 399
rect 1428 405 1440 411
rect 1524 417 1536 420
rect 1524 411 1527 417
rect 1533 411 1536 417
rect 1428 399 1431 405
rect 1437 399 1440 405
rect 1428 396 1440 399
rect 1452 405 1512 408
rect 1452 399 1455 405
rect 1461 399 1503 405
rect 1509 399 1512 405
rect 1452 396 1512 399
rect 1524 405 1536 411
rect 1524 399 1527 405
rect 1533 399 1536 405
rect 1524 396 1536 399
rect 1572 429 1584 471
rect 1596 453 1608 456
rect 1596 447 1599 453
rect 1605 447 1608 453
rect 1596 444 1608 447
rect 1572 423 1575 429
rect 1581 423 1584 429
rect 1572 417 1584 423
rect 1572 411 1575 417
rect 1581 411 1584 417
rect 1572 405 1584 411
rect 1572 399 1575 405
rect 1581 399 1584 405
rect 1572 396 1584 399
rect 12 381 24 384
rect 12 375 15 381
rect 21 375 24 381
rect 12 372 24 375
rect -60 333 -48 336
rect -60 327 -57 333
rect -51 327 -48 333
rect -60 285 -48 327
rect -60 279 -57 285
rect -51 279 -48 285
rect -60 237 -48 279
rect -60 231 -57 237
rect -51 231 -48 237
rect -60 189 -48 231
rect -60 183 -57 189
rect -51 183 -48 189
rect -60 93 -48 183
rect -60 87 -57 93
rect -51 87 -48 93
rect -60 45 -48 87
rect -60 39 -57 45
rect -51 39 -48 45
rect -60 33 -48 39
rect -60 27 -57 33
rect -51 27 -48 33
rect -60 21 -48 27
rect -60 15 -57 21
rect -51 15 -48 21
rect -60 -3 -48 15
rect -60 -9 -57 -3
rect -51 -9 -48 -3
rect -60 -12 -48 -9
rect -12 333 0 336
rect -12 327 -9 333
rect -3 327 0 333
rect -12 285 0 327
rect -12 279 -9 285
rect -3 279 0 285
rect -12 237 0 279
rect -12 231 -9 237
rect -3 231 0 237
rect -12 189 0 231
rect -12 183 -9 189
rect -3 183 0 189
rect -12 93 0 183
rect -12 87 -9 93
rect -3 87 0 93
rect -12 45 0 87
rect 36 165 48 396
rect 60 381 72 384
rect 60 375 63 381
rect 69 375 72 381
rect 60 372 72 375
rect 108 381 120 384
rect 108 375 111 381
rect 117 375 120 381
rect 108 372 120 375
rect 36 159 39 165
rect 45 159 48 165
rect 36 117 48 159
rect 36 111 39 117
rect 45 111 48 117
rect 12 69 24 72
rect 12 63 15 69
rect 21 63 24 69
rect 12 60 24 63
rect -12 39 -9 45
rect -3 39 0 45
rect -12 33 0 39
rect -12 27 -9 33
rect -3 27 0 33
rect -12 21 0 27
rect -12 15 -9 21
rect -3 15 0 21
rect -12 -3 0 15
rect 36 45 48 111
rect 132 165 144 396
rect 156 381 168 384
rect 156 375 159 381
rect 165 375 168 381
rect 156 372 168 375
rect 204 381 216 384
rect 204 375 207 381
rect 213 375 216 381
rect 204 372 216 375
rect 252 381 264 384
rect 252 375 255 381
rect 261 375 264 381
rect 252 372 264 375
rect 132 159 135 165
rect 141 159 144 165
rect 132 117 144 159
rect 132 111 135 117
rect 141 111 144 117
rect 60 69 72 72
rect 60 63 63 69
rect 69 63 72 69
rect 60 60 72 63
rect 108 69 120 72
rect 108 63 111 69
rect 117 63 120 69
rect 108 60 120 63
rect 36 39 39 45
rect 45 39 48 45
rect 36 33 48 39
rect 36 27 39 33
rect 45 27 48 33
rect 36 21 48 27
rect 36 15 39 21
rect 45 15 48 21
rect 36 12 48 15
rect 84 45 96 48
rect 84 39 87 45
rect 93 39 96 45
rect 84 33 96 39
rect 84 27 87 33
rect 93 27 96 33
rect 84 21 96 27
rect 84 15 87 21
rect 93 15 96 21
rect 84 12 96 15
rect 132 45 144 111
rect 180 333 192 336
rect 180 327 183 333
rect 189 327 192 333
rect 180 285 192 327
rect 180 279 183 285
rect 189 279 192 285
rect 180 237 192 279
rect 180 231 183 237
rect 189 231 192 237
rect 180 189 192 231
rect 180 183 183 189
rect 189 183 192 189
rect 180 93 192 183
rect 180 87 183 93
rect 189 87 192 93
rect 156 69 168 72
rect 156 63 159 69
rect 165 63 168 69
rect 156 60 168 63
rect 132 39 135 45
rect 141 39 144 45
rect 132 33 144 39
rect 132 27 135 33
rect 141 27 144 33
rect 132 21 144 27
rect 132 15 135 21
rect 141 15 144 21
rect 132 12 144 15
rect 180 45 192 87
rect 276 141 288 396
rect 300 381 312 384
rect 300 375 303 381
rect 309 375 312 381
rect 300 372 312 375
rect 348 381 360 384
rect 348 375 351 381
rect 357 375 360 381
rect 348 372 360 375
rect 396 381 408 384
rect 396 375 399 381
rect 405 375 408 381
rect 396 372 408 375
rect 444 381 456 384
rect 444 375 447 381
rect 453 375 456 381
rect 444 372 456 375
rect 276 135 279 141
rect 285 135 288 141
rect 204 69 216 72
rect 204 63 207 69
rect 213 63 216 69
rect 204 60 216 63
rect 252 69 264 72
rect 252 63 255 69
rect 261 63 264 69
rect 252 60 264 63
rect 180 39 183 45
rect 189 39 192 45
rect 180 33 192 39
rect 180 27 183 33
rect 189 27 192 33
rect 180 21 192 27
rect 180 15 183 21
rect 189 15 192 21
rect -12 -9 -9 -3
rect -3 -9 0 -3
rect -12 -12 0 -9
rect 180 -3 192 15
rect 276 45 288 135
rect 372 333 384 336
rect 372 327 375 333
rect 381 327 384 333
rect 372 285 384 327
rect 372 279 375 285
rect 381 279 384 285
rect 372 237 384 279
rect 372 231 375 237
rect 381 231 384 237
rect 372 189 384 231
rect 372 183 375 189
rect 381 183 384 189
rect 372 93 384 183
rect 372 87 375 93
rect 381 87 384 93
rect 300 69 312 72
rect 300 63 303 69
rect 309 63 312 69
rect 300 60 312 63
rect 348 69 360 72
rect 348 63 351 69
rect 357 63 360 69
rect 348 60 360 63
rect 276 39 279 45
rect 285 39 288 45
rect 276 33 288 39
rect 276 27 279 33
rect 285 27 288 33
rect 276 21 288 27
rect 276 15 279 21
rect 285 15 288 21
rect 276 12 288 15
rect 372 45 384 87
rect 468 261 480 396
rect 492 381 504 384
rect 492 375 495 381
rect 501 375 504 381
rect 492 372 504 375
rect 540 381 552 384
rect 540 375 543 381
rect 549 375 552 381
rect 540 372 552 375
rect 588 381 600 384
rect 588 375 591 381
rect 597 375 600 381
rect 588 372 600 375
rect 468 255 471 261
rect 477 255 480 261
rect 396 69 408 72
rect 396 63 399 69
rect 405 63 408 69
rect 396 60 408 63
rect 444 69 456 72
rect 444 63 447 69
rect 453 63 456 69
rect 444 60 456 63
rect 372 39 375 45
rect 381 39 384 45
rect 372 33 384 39
rect 372 27 375 33
rect 381 27 384 33
rect 372 21 384 27
rect 372 15 375 21
rect 381 15 384 21
rect 180 -9 183 -3
rect 189 -9 192 -3
rect 180 -12 192 -9
rect 372 -3 384 15
rect 468 45 480 255
rect 564 333 576 336
rect 564 327 567 333
rect 573 327 576 333
rect 564 285 576 327
rect 564 279 567 285
rect 573 279 576 285
rect 564 237 576 279
rect 564 231 567 237
rect 573 231 576 237
rect 564 189 576 231
rect 564 183 567 189
rect 573 183 576 189
rect 564 93 576 183
rect 564 87 567 93
rect 573 87 576 93
rect 492 69 504 72
rect 492 63 495 69
rect 501 63 504 69
rect 492 60 504 63
rect 540 69 552 72
rect 540 63 543 69
rect 549 63 552 69
rect 540 60 552 63
rect 468 39 471 45
rect 477 39 480 45
rect 468 33 480 39
rect 468 27 471 33
rect 477 27 480 33
rect 468 21 480 27
rect 468 15 471 21
rect 477 15 480 21
rect 468 12 480 15
rect 564 45 576 87
rect 612 165 624 396
rect 636 381 648 384
rect 636 375 639 381
rect 645 375 648 381
rect 636 372 648 375
rect 684 381 696 384
rect 684 375 687 381
rect 693 375 696 381
rect 684 372 696 375
rect 612 159 615 165
rect 621 159 624 165
rect 612 117 624 159
rect 612 111 615 117
rect 621 111 624 117
rect 588 69 600 72
rect 588 63 591 69
rect 597 63 600 69
rect 588 60 600 63
rect 564 39 567 45
rect 573 39 576 45
rect 564 33 576 39
rect 564 27 567 33
rect 573 27 576 33
rect 564 21 576 27
rect 564 15 567 21
rect 573 15 576 21
rect 372 -9 375 -3
rect 381 -9 384 -3
rect 372 -12 384 -9
rect 564 -3 576 15
rect 612 45 624 111
rect 708 165 720 396
rect 732 381 744 384
rect 732 375 735 381
rect 741 375 744 381
rect 732 372 744 375
rect 780 381 792 384
rect 780 375 783 381
rect 789 375 792 381
rect 780 372 792 375
rect 708 159 711 165
rect 717 159 720 165
rect 708 117 720 159
rect 708 111 711 117
rect 717 111 720 117
rect 636 69 648 72
rect 636 63 639 69
rect 645 63 648 69
rect 636 60 648 63
rect 684 69 696 72
rect 684 63 687 69
rect 693 63 696 69
rect 684 60 696 63
rect 612 39 615 45
rect 621 39 624 45
rect 612 33 624 39
rect 612 27 615 33
rect 621 27 624 33
rect 612 21 624 27
rect 612 15 615 21
rect 621 15 624 21
rect 612 12 624 15
rect 660 45 672 48
rect 660 39 663 45
rect 669 39 672 45
rect 660 33 672 39
rect 660 27 663 33
rect 669 27 672 33
rect 660 21 672 27
rect 660 15 663 21
rect 669 15 672 21
rect 660 12 672 15
rect 708 45 720 111
rect 756 333 768 336
rect 756 327 759 333
rect 765 327 768 333
rect 756 285 768 327
rect 756 279 759 285
rect 765 279 768 285
rect 756 237 768 279
rect 756 231 759 237
rect 765 231 768 237
rect 756 189 768 231
rect 756 183 759 189
rect 765 183 768 189
rect 756 93 768 183
rect 756 87 759 93
rect 765 87 768 93
rect 732 69 744 72
rect 732 63 735 69
rect 741 63 744 69
rect 732 60 744 63
rect 708 39 711 45
rect 717 39 720 45
rect 708 33 720 39
rect 708 27 711 33
rect 717 27 720 33
rect 708 21 720 27
rect 708 15 711 21
rect 717 15 720 21
rect 708 12 720 15
rect 756 45 768 87
rect 804 165 816 396
rect 828 381 840 384
rect 828 375 831 381
rect 837 375 840 381
rect 828 372 840 375
rect 876 381 888 384
rect 876 375 879 381
rect 885 375 888 381
rect 876 372 888 375
rect 804 159 807 165
rect 813 159 816 165
rect 804 117 816 159
rect 804 111 807 117
rect 813 111 816 117
rect 780 69 792 72
rect 780 63 783 69
rect 789 63 792 69
rect 780 60 792 63
rect 756 39 759 45
rect 765 39 768 45
rect 756 33 768 39
rect 756 27 759 33
rect 765 27 768 33
rect 756 21 768 27
rect 756 15 759 21
rect 765 15 768 21
rect 564 -9 567 -3
rect 573 -9 576 -3
rect 564 -12 576 -9
rect 756 -3 768 15
rect 804 45 816 111
rect 900 165 912 396
rect 924 381 936 384
rect 924 375 927 381
rect 933 375 936 381
rect 924 372 936 375
rect 972 381 984 384
rect 972 375 975 381
rect 981 375 984 381
rect 972 372 984 375
rect 1020 381 1032 384
rect 1020 375 1023 381
rect 1029 375 1032 381
rect 1020 372 1032 375
rect 900 159 903 165
rect 909 159 912 165
rect 900 117 912 159
rect 900 111 903 117
rect 909 111 912 117
rect 828 69 840 72
rect 828 63 831 69
rect 837 63 840 69
rect 828 60 840 63
rect 876 69 888 72
rect 876 63 879 69
rect 885 63 888 69
rect 876 60 888 63
rect 804 39 807 45
rect 813 39 816 45
rect 804 33 816 39
rect 804 27 807 33
rect 813 27 816 33
rect 804 21 816 27
rect 804 15 807 21
rect 813 15 816 21
rect 804 12 816 15
rect 852 45 864 48
rect 852 39 855 45
rect 861 39 864 45
rect 852 33 864 39
rect 852 27 855 33
rect 861 27 864 33
rect 852 21 864 27
rect 852 15 855 21
rect 861 15 864 21
rect 852 12 864 15
rect 900 45 912 111
rect 948 333 960 336
rect 948 327 951 333
rect 957 327 960 333
rect 948 285 960 327
rect 948 279 951 285
rect 957 279 960 285
rect 948 237 960 279
rect 948 231 951 237
rect 957 231 960 237
rect 948 189 960 231
rect 948 183 951 189
rect 957 183 960 189
rect 948 93 960 183
rect 948 87 951 93
rect 957 87 960 93
rect 924 69 936 72
rect 924 63 927 69
rect 933 63 936 69
rect 924 60 936 63
rect 900 39 903 45
rect 909 39 912 45
rect 900 33 912 39
rect 900 27 903 33
rect 909 27 912 33
rect 900 21 912 27
rect 900 15 903 21
rect 909 15 912 21
rect 900 12 912 15
rect 948 45 960 87
rect 1044 261 1056 396
rect 1068 381 1080 384
rect 1068 375 1071 381
rect 1077 375 1080 381
rect 1068 372 1080 375
rect 1116 381 1128 384
rect 1116 375 1119 381
rect 1125 375 1128 381
rect 1116 372 1128 375
rect 1164 381 1176 384
rect 1164 375 1167 381
rect 1173 375 1176 381
rect 1164 372 1176 375
rect 1212 381 1224 384
rect 1212 375 1215 381
rect 1221 375 1224 381
rect 1212 372 1224 375
rect 1044 255 1047 261
rect 1053 255 1056 261
rect 972 69 984 72
rect 972 63 975 69
rect 981 63 984 69
rect 972 60 984 63
rect 1020 69 1032 72
rect 1020 63 1023 69
rect 1029 63 1032 69
rect 1020 60 1032 63
rect 948 39 951 45
rect 957 39 960 45
rect 948 33 960 39
rect 948 27 951 33
rect 957 27 960 33
rect 948 21 960 27
rect 948 15 951 21
rect 957 15 960 21
rect 756 -9 759 -3
rect 765 -9 768 -3
rect 756 -12 768 -9
rect 948 -3 960 15
rect 1044 45 1056 255
rect 1140 333 1152 336
rect 1140 327 1143 333
rect 1149 327 1152 333
rect 1140 285 1152 327
rect 1140 279 1143 285
rect 1149 279 1152 285
rect 1140 237 1152 279
rect 1140 231 1143 237
rect 1149 231 1152 237
rect 1140 189 1152 231
rect 1140 183 1143 189
rect 1149 183 1152 189
rect 1140 93 1152 183
rect 1140 87 1143 93
rect 1149 87 1152 93
rect 1068 69 1080 72
rect 1068 63 1071 69
rect 1077 63 1080 69
rect 1068 60 1080 63
rect 1116 69 1128 72
rect 1116 63 1119 69
rect 1125 63 1128 69
rect 1116 60 1128 63
rect 1044 39 1047 45
rect 1053 39 1056 45
rect 1044 33 1056 39
rect 1044 27 1047 33
rect 1053 27 1056 33
rect 1044 21 1056 27
rect 1044 15 1047 21
rect 1053 15 1056 21
rect 1044 12 1056 15
rect 1140 45 1152 87
rect 1236 141 1248 396
rect 1260 381 1272 384
rect 1260 375 1263 381
rect 1269 375 1272 381
rect 1260 372 1272 375
rect 1308 381 1320 384
rect 1308 375 1311 381
rect 1317 375 1320 381
rect 1308 372 1320 375
rect 1356 381 1368 384
rect 1356 375 1359 381
rect 1365 375 1368 381
rect 1356 372 1368 375
rect 1236 135 1239 141
rect 1245 135 1248 141
rect 1164 69 1176 72
rect 1164 63 1167 69
rect 1173 63 1176 69
rect 1164 60 1176 63
rect 1212 69 1224 72
rect 1212 63 1215 69
rect 1221 63 1224 69
rect 1212 60 1224 63
rect 1140 39 1143 45
rect 1149 39 1152 45
rect 1140 33 1152 39
rect 1140 27 1143 33
rect 1149 27 1152 33
rect 1140 21 1152 27
rect 1140 15 1143 21
rect 1149 15 1152 21
rect 948 -9 951 -3
rect 957 -9 960 -3
rect 948 -12 960 -9
rect 1140 -3 1152 15
rect 1236 45 1248 135
rect 1332 333 1344 336
rect 1332 327 1335 333
rect 1341 327 1344 333
rect 1332 285 1344 327
rect 1380 324 1392 396
rect 1404 381 1416 384
rect 1404 375 1407 381
rect 1413 375 1416 381
rect 1404 372 1416 375
rect 1452 381 1464 384
rect 1452 375 1455 381
rect 1461 375 1464 381
rect 1452 372 1464 375
rect 1332 279 1335 285
rect 1341 279 1344 285
rect 1332 237 1344 279
rect 1332 231 1335 237
rect 1341 231 1344 237
rect 1332 189 1344 231
rect 1332 183 1335 189
rect 1341 183 1344 189
rect 1332 93 1344 183
rect 1332 87 1335 93
rect 1341 87 1344 93
rect 1260 69 1272 72
rect 1260 63 1263 69
rect 1269 63 1272 69
rect 1260 60 1272 63
rect 1308 69 1320 72
rect 1308 63 1311 69
rect 1317 63 1320 69
rect 1308 60 1320 63
rect 1236 39 1239 45
rect 1245 39 1248 45
rect 1236 33 1248 39
rect 1236 27 1239 33
rect 1245 27 1248 33
rect 1236 21 1248 27
rect 1236 15 1239 21
rect 1245 15 1248 21
rect 1236 12 1248 15
rect 1332 45 1344 87
rect 1380 165 1392 312
rect 1380 159 1383 165
rect 1389 159 1392 165
rect 1380 117 1392 159
rect 1380 111 1383 117
rect 1389 111 1392 117
rect 1356 69 1368 72
rect 1356 63 1359 69
rect 1365 63 1368 69
rect 1356 60 1368 63
rect 1332 39 1335 45
rect 1341 39 1344 45
rect 1332 33 1344 39
rect 1332 27 1335 33
rect 1341 27 1344 33
rect 1332 21 1344 27
rect 1332 15 1335 21
rect 1341 15 1344 21
rect 1140 -9 1143 -3
rect 1149 -9 1152 -3
rect 1140 -12 1152 -9
rect 1332 -3 1344 15
rect 1380 45 1392 111
rect 1476 165 1488 396
rect 1500 381 1512 384
rect 1500 375 1503 381
rect 1509 375 1512 381
rect 1500 372 1512 375
rect 1476 159 1479 165
rect 1485 159 1488 165
rect 1476 117 1488 159
rect 1476 111 1479 117
rect 1485 111 1488 117
rect 1404 69 1416 72
rect 1404 63 1407 69
rect 1413 63 1416 69
rect 1404 60 1416 63
rect 1452 69 1464 72
rect 1452 63 1455 69
rect 1461 63 1464 69
rect 1452 60 1464 63
rect 1380 39 1383 45
rect 1389 39 1392 45
rect 1380 33 1392 39
rect 1380 27 1383 33
rect 1389 27 1392 33
rect 1380 21 1392 27
rect 1380 15 1383 21
rect 1389 15 1392 21
rect 1380 12 1392 15
rect 1428 45 1440 48
rect 1428 39 1431 45
rect 1437 39 1440 45
rect 1428 33 1440 39
rect 1428 27 1431 33
rect 1437 27 1440 33
rect 1428 21 1440 27
rect 1428 15 1431 21
rect 1437 15 1440 21
rect 1428 12 1440 15
rect 1476 45 1488 111
rect 1524 333 1536 336
rect 1524 327 1527 333
rect 1533 327 1536 333
rect 1524 285 1536 327
rect 1524 279 1527 285
rect 1533 279 1536 285
rect 1524 237 1536 279
rect 1524 231 1527 237
rect 1533 231 1536 237
rect 1524 189 1536 231
rect 1524 183 1527 189
rect 1533 183 1536 189
rect 1524 93 1536 183
rect 1524 87 1527 93
rect 1533 87 1536 93
rect 1500 69 1512 72
rect 1500 63 1503 69
rect 1509 63 1512 69
rect 1500 60 1512 63
rect 1476 39 1479 45
rect 1485 39 1488 45
rect 1476 33 1488 39
rect 1476 27 1479 33
rect 1485 27 1488 33
rect 1476 21 1488 27
rect 1476 15 1479 21
rect 1485 15 1488 21
rect 1476 12 1488 15
rect 1524 45 1536 87
rect 1524 39 1527 45
rect 1533 39 1536 45
rect 1524 33 1536 39
rect 1524 27 1527 33
rect 1533 27 1536 33
rect 1524 21 1536 27
rect 1524 15 1527 21
rect 1533 15 1536 21
rect 1332 -9 1335 -3
rect 1341 -9 1344 -3
rect 1332 -12 1344 -9
rect 1524 -3 1536 15
rect 1524 -9 1527 -3
rect 1533 -9 1536 -3
rect 1524 -12 1536 -9
rect 1572 333 1584 336
rect 1572 327 1575 333
rect 1581 327 1584 333
rect 1572 285 1584 327
rect 1572 279 1575 285
rect 1581 279 1584 285
rect 1572 237 1584 279
rect 1572 231 1575 237
rect 1581 231 1584 237
rect 1572 189 1584 231
rect 1572 183 1575 189
rect 1581 183 1584 189
rect 1572 93 1584 183
rect 1572 87 1575 93
rect 1581 87 1584 93
rect 1572 45 1584 87
rect 1572 39 1575 45
rect 1581 39 1584 45
rect 1572 33 1584 39
rect 1572 27 1575 33
rect 1581 27 1584 33
rect 1572 21 1584 27
rect 1572 15 1575 21
rect 1581 15 1584 21
rect 1572 -3 1584 15
rect 1572 -9 1575 -3
rect 1581 -9 1584 -3
rect 1572 -12 1584 -9
<< via2 >>
rect -81 591 -75 597
rect 1599 591 1605 597
rect -33 567 -27 573
rect 15 567 21 573
rect 63 567 69 573
rect 111 567 117 573
rect 159 567 165 573
rect 207 567 213 573
rect 255 567 261 573
rect 303 567 309 573
rect 351 567 357 573
rect 399 567 405 573
rect 447 567 453 573
rect 495 567 501 573
rect 543 567 549 573
rect 591 567 597 573
rect 639 567 645 573
rect 687 567 693 573
rect 735 567 741 573
rect 783 567 789 573
rect 831 567 837 573
rect 879 567 885 573
rect 927 567 933 573
rect 975 567 981 573
rect 1023 567 1029 573
rect 1071 567 1077 573
rect 1119 567 1125 573
rect 1167 567 1173 573
rect 1215 567 1221 573
rect 1263 567 1269 573
rect 1311 567 1317 573
rect 1359 567 1365 573
rect 1407 567 1413 573
rect 1455 567 1461 573
rect 1503 567 1509 573
rect 1551 567 1557 573
rect -81 543 -75 549
rect -81 531 -75 537
rect -81 519 -75 525
rect -57 471 -51 477
rect -81 447 -75 453
rect 15 543 21 549
rect 15 531 21 537
rect 15 519 21 525
rect -9 471 -3 477
rect -33 447 -27 453
rect -57 423 -51 429
rect -57 411 -51 417
rect -57 399 -51 405
rect 63 543 69 549
rect 63 531 69 537
rect 63 519 69 525
rect 39 471 45 477
rect 15 447 21 453
rect 111 543 117 549
rect 111 531 117 537
rect 111 519 117 525
rect 87 471 93 477
rect 63 447 69 453
rect 159 543 165 549
rect 159 531 165 537
rect 159 519 165 525
rect 135 471 141 477
rect 111 447 117 453
rect 207 543 213 549
rect 207 531 213 537
rect 207 519 213 525
rect 183 471 189 477
rect 159 447 165 453
rect 255 543 261 549
rect 255 531 261 537
rect 255 519 261 525
rect 231 471 237 477
rect 207 447 213 453
rect 303 543 309 549
rect 303 531 309 537
rect 303 519 309 525
rect 279 471 285 477
rect 255 447 261 453
rect 351 543 357 549
rect 351 531 357 537
rect 351 519 357 525
rect 327 471 333 477
rect 303 447 309 453
rect 399 543 405 549
rect 399 531 405 537
rect 399 519 405 525
rect 375 471 381 477
rect 351 447 357 453
rect 447 543 453 549
rect 447 531 453 537
rect 447 519 453 525
rect 423 471 429 477
rect 399 447 405 453
rect 495 543 501 549
rect 495 531 501 537
rect 495 519 501 525
rect 471 471 477 477
rect 447 447 453 453
rect 543 543 549 549
rect 543 531 549 537
rect 543 519 549 525
rect 519 471 525 477
rect 495 447 501 453
rect 591 543 597 549
rect 591 531 597 537
rect 591 519 597 525
rect 567 471 573 477
rect 543 447 549 453
rect 639 543 645 549
rect 639 531 645 537
rect 639 519 645 525
rect 615 471 621 477
rect 591 447 597 453
rect 687 543 693 549
rect 687 531 693 537
rect 687 519 693 525
rect 663 471 669 477
rect 639 447 645 453
rect 735 543 741 549
rect 735 531 741 537
rect 735 519 741 525
rect 711 471 717 477
rect 687 447 693 453
rect 783 543 789 549
rect 783 531 789 537
rect 783 519 789 525
rect 759 471 765 477
rect 735 447 741 453
rect 831 543 837 549
rect 831 531 837 537
rect 831 519 837 525
rect 807 471 813 477
rect 783 447 789 453
rect 879 543 885 549
rect 879 531 885 537
rect 879 519 885 525
rect 855 471 861 477
rect 831 447 837 453
rect 927 543 933 549
rect 927 531 933 537
rect 927 519 933 525
rect 903 471 909 477
rect 879 447 885 453
rect 975 543 981 549
rect 975 531 981 537
rect 975 519 981 525
rect 951 471 957 477
rect 927 447 933 453
rect 1023 543 1029 549
rect 1023 531 1029 537
rect 1023 519 1029 525
rect 999 471 1005 477
rect 975 447 981 453
rect 1071 543 1077 549
rect 1071 531 1077 537
rect 1071 519 1077 525
rect 1047 471 1053 477
rect 1023 447 1029 453
rect 1119 543 1125 549
rect 1119 531 1125 537
rect 1119 519 1125 525
rect 1095 471 1101 477
rect 1071 447 1077 453
rect 1167 543 1173 549
rect 1167 531 1173 537
rect 1167 519 1173 525
rect 1143 471 1149 477
rect 1119 447 1125 453
rect 1215 543 1221 549
rect 1215 531 1221 537
rect 1215 519 1221 525
rect 1191 471 1197 477
rect 1167 447 1173 453
rect 1263 543 1269 549
rect 1263 531 1269 537
rect 1263 519 1269 525
rect 1239 471 1245 477
rect 1215 447 1221 453
rect 1311 543 1317 549
rect 1311 531 1317 537
rect 1311 519 1317 525
rect 1287 471 1293 477
rect 1263 447 1269 453
rect 1359 543 1365 549
rect 1359 531 1365 537
rect 1359 519 1365 525
rect 1335 471 1341 477
rect 1311 447 1317 453
rect 1407 543 1413 549
rect 1407 531 1413 537
rect 1407 519 1413 525
rect 1383 471 1389 477
rect 1359 447 1365 453
rect 1455 543 1461 549
rect 1455 531 1461 537
rect 1455 519 1461 525
rect 1431 471 1437 477
rect 1407 447 1413 453
rect 1503 543 1509 549
rect 1503 531 1509 537
rect 1503 519 1509 525
rect 1479 471 1485 477
rect 1455 447 1461 453
rect 1527 471 1533 477
rect 1503 447 1509 453
rect 1599 543 1605 549
rect 1599 531 1605 537
rect 1599 519 1605 525
rect 1575 471 1581 477
rect 1551 447 1557 453
rect -9 423 -3 429
rect 39 423 45 429
rect 87 423 93 429
rect 183 423 189 429
rect 279 423 285 429
rect 375 423 381 429
rect 471 423 477 429
rect 567 423 573 429
rect 615 423 621 429
rect 663 423 669 429
rect 759 423 765 429
rect 855 423 861 429
rect 903 423 909 429
rect 951 423 957 429
rect 1047 423 1053 429
rect 1143 423 1149 429
rect 1239 423 1245 429
rect 1335 423 1341 429
rect 1431 423 1437 429
rect 1479 423 1485 429
rect 1527 423 1533 429
rect -9 411 -3 417
rect 87 411 93 417
rect -9 399 -3 405
rect 183 411 189 417
rect 87 399 93 405
rect 375 411 381 417
rect 183 399 189 405
rect 567 411 573 417
rect 375 399 381 405
rect 663 411 669 417
rect 567 399 573 405
rect 759 411 765 417
rect 663 399 669 405
rect 855 411 861 417
rect 759 399 765 405
rect 951 411 957 417
rect 855 399 861 405
rect 1143 411 1149 417
rect 951 399 957 405
rect 1335 411 1341 417
rect 1143 399 1149 405
rect 1431 411 1437 417
rect 1335 399 1341 405
rect 1527 411 1533 417
rect 1431 399 1437 405
rect 1527 399 1533 405
rect 1599 447 1605 453
rect 1575 423 1581 429
rect 1575 411 1581 417
rect 1575 399 1581 405
rect 15 375 21 381
rect -57 327 -51 333
rect -57 279 -51 285
rect -57 231 -51 237
rect -57 183 -51 189
rect -57 87 -51 93
rect -57 39 -51 45
rect -57 27 -51 33
rect -57 15 -51 21
rect -9 327 -3 333
rect -9 279 -3 285
rect -9 231 -3 237
rect -9 183 -3 189
rect -9 87 -3 93
rect 63 375 69 381
rect 111 375 117 381
rect 39 159 45 165
rect 39 111 45 117
rect 15 63 21 69
rect -9 39 -3 45
rect -9 27 -3 33
rect -9 15 -3 21
rect 159 375 165 381
rect 207 375 213 381
rect 255 375 261 381
rect 135 159 141 165
rect 135 111 141 117
rect 63 63 69 69
rect 111 63 117 69
rect 87 39 93 45
rect 87 27 93 33
rect 87 15 93 21
rect 183 327 189 333
rect 183 279 189 285
rect 183 231 189 237
rect 183 183 189 189
rect 183 87 189 93
rect 159 63 165 69
rect 303 375 309 381
rect 351 375 357 381
rect 399 375 405 381
rect 447 375 453 381
rect 279 135 285 141
rect 207 63 213 69
rect 255 63 261 69
rect 183 39 189 45
rect 183 27 189 33
rect 183 15 189 21
rect 375 327 381 333
rect 375 279 381 285
rect 375 231 381 237
rect 375 183 381 189
rect 375 87 381 93
rect 303 63 309 69
rect 351 63 357 69
rect 495 375 501 381
rect 543 375 549 381
rect 591 375 597 381
rect 471 255 477 261
rect 399 63 405 69
rect 447 63 453 69
rect 375 39 381 45
rect 375 27 381 33
rect 375 15 381 21
rect 567 327 573 333
rect 567 279 573 285
rect 567 231 573 237
rect 567 183 573 189
rect 567 87 573 93
rect 495 63 501 69
rect 543 63 549 69
rect 639 375 645 381
rect 687 375 693 381
rect 615 159 621 165
rect 615 111 621 117
rect 591 63 597 69
rect 567 39 573 45
rect 567 27 573 33
rect 567 15 573 21
rect 735 375 741 381
rect 783 375 789 381
rect 711 159 717 165
rect 711 111 717 117
rect 639 63 645 69
rect 687 63 693 69
rect 663 39 669 45
rect 663 27 669 33
rect 663 15 669 21
rect 759 327 765 333
rect 759 279 765 285
rect 759 231 765 237
rect 759 183 765 189
rect 759 87 765 93
rect 735 63 741 69
rect 831 375 837 381
rect 879 375 885 381
rect 807 159 813 165
rect 807 111 813 117
rect 783 63 789 69
rect 759 39 765 45
rect 759 27 765 33
rect 759 15 765 21
rect 927 375 933 381
rect 975 375 981 381
rect 1023 375 1029 381
rect 903 159 909 165
rect 903 111 909 117
rect 831 63 837 69
rect 879 63 885 69
rect 855 39 861 45
rect 855 27 861 33
rect 855 15 861 21
rect 951 327 957 333
rect 951 279 957 285
rect 951 231 957 237
rect 951 183 957 189
rect 951 87 957 93
rect 927 63 933 69
rect 1071 375 1077 381
rect 1119 375 1125 381
rect 1167 375 1173 381
rect 1215 375 1221 381
rect 1047 255 1053 261
rect 975 63 981 69
rect 1023 63 1029 69
rect 951 39 957 45
rect 951 27 957 33
rect 951 15 957 21
rect 1143 327 1149 333
rect 1143 279 1149 285
rect 1143 231 1149 237
rect 1143 183 1149 189
rect 1143 87 1149 93
rect 1071 63 1077 69
rect 1119 63 1125 69
rect 1263 375 1269 381
rect 1311 375 1317 381
rect 1359 375 1365 381
rect 1239 135 1245 141
rect 1167 63 1173 69
rect 1215 63 1221 69
rect 1143 39 1149 45
rect 1143 27 1149 33
rect 1143 15 1149 21
rect 1335 327 1341 333
rect 1407 375 1413 381
rect 1455 375 1461 381
rect 1335 279 1341 285
rect 1335 231 1341 237
rect 1335 183 1341 189
rect 1335 87 1341 93
rect 1263 63 1269 69
rect 1311 63 1317 69
rect 1383 159 1389 165
rect 1383 111 1389 117
rect 1359 63 1365 69
rect 1335 39 1341 45
rect 1335 27 1341 33
rect 1335 15 1341 21
rect 1503 375 1509 381
rect 1479 159 1485 165
rect 1479 111 1485 117
rect 1407 63 1413 69
rect 1455 63 1461 69
rect 1431 39 1437 45
rect 1431 27 1437 33
rect 1431 15 1437 21
rect 1527 327 1533 333
rect 1527 279 1533 285
rect 1527 231 1533 237
rect 1527 183 1533 189
rect 1527 87 1533 93
rect 1503 63 1509 69
rect 1527 39 1533 45
rect 1527 27 1533 33
rect 1527 15 1533 21
rect 1575 327 1581 333
rect 1575 279 1581 285
rect 1575 231 1581 237
rect 1575 183 1581 189
rect 1575 87 1581 93
rect 1575 39 1581 45
rect 1575 27 1581 33
rect 1575 15 1581 21
<< mimcap >>
rect -48 -72 1572 -60
rect -48 -156 -36 -72
rect 1560 -156 1572 -72
rect -48 -168 1572 -156
<< mimcapcontact >>
rect -36 -156 1560 -72
<< metal3 >>
rect -108 597 1632 600
rect -108 591 -81 597
rect -75 591 1599 597
rect 1605 591 1632 597
rect -108 582 1632 591
rect -108 573 1632 576
rect -108 567 -33 573
rect -27 567 15 573
rect 21 567 63 573
rect 69 567 111 573
rect 117 567 159 573
rect 165 567 207 573
rect 213 567 255 573
rect 261 567 303 573
rect 309 567 351 573
rect 357 567 399 573
rect 405 567 447 573
rect 453 567 495 573
rect 501 567 543 573
rect 549 567 591 573
rect 597 567 639 573
rect 645 567 687 573
rect 693 567 735 573
rect 741 567 783 573
rect 789 567 831 573
rect 837 567 879 573
rect 885 567 927 573
rect 933 567 975 573
rect 981 567 1023 573
rect 1029 567 1071 573
rect 1077 567 1119 573
rect 1125 567 1167 573
rect 1173 567 1215 573
rect 1221 567 1263 573
rect 1269 567 1311 573
rect 1317 567 1359 573
rect 1365 567 1407 573
rect 1413 567 1455 573
rect 1461 567 1503 573
rect 1509 567 1551 573
rect 1557 567 1632 573
rect -108 564 1632 567
rect -108 549 1632 558
rect -108 543 -81 549
rect -75 543 15 549
rect 21 543 63 549
rect 69 543 111 549
rect 117 543 159 549
rect 165 543 207 549
rect 213 543 255 549
rect 261 543 303 549
rect 309 543 351 549
rect 357 543 399 549
rect 405 543 447 549
rect 453 543 495 549
rect 501 543 543 549
rect 549 543 591 549
rect 597 543 639 549
rect 645 543 687 549
rect 693 543 735 549
rect 741 543 783 549
rect 789 543 831 549
rect 837 543 879 549
rect 885 543 927 549
rect 933 543 975 549
rect 981 543 1023 549
rect 1029 543 1071 549
rect 1077 543 1119 549
rect 1125 543 1167 549
rect 1173 543 1215 549
rect 1221 543 1263 549
rect 1269 543 1311 549
rect 1317 543 1359 549
rect 1365 543 1407 549
rect 1413 543 1455 549
rect 1461 543 1503 549
rect 1509 543 1599 549
rect 1605 543 1632 549
rect -108 537 1632 543
rect -108 531 -81 537
rect -75 531 15 537
rect 21 531 63 537
rect 69 531 111 537
rect 117 531 159 537
rect 165 531 207 537
rect 213 531 255 537
rect 261 531 303 537
rect 309 531 351 537
rect 357 531 399 537
rect 405 531 447 537
rect 453 531 495 537
rect 501 531 543 537
rect 549 531 591 537
rect 597 531 639 537
rect 645 531 687 537
rect 693 531 735 537
rect 741 531 783 537
rect 789 531 831 537
rect 837 531 879 537
rect 885 531 927 537
rect 933 531 975 537
rect 981 531 1023 537
rect 1029 531 1071 537
rect 1077 531 1119 537
rect 1125 531 1167 537
rect 1173 531 1215 537
rect 1221 531 1263 537
rect 1269 531 1311 537
rect 1317 531 1359 537
rect 1365 531 1407 537
rect 1413 531 1455 537
rect 1461 531 1503 537
rect 1509 531 1599 537
rect 1605 531 1632 537
rect -108 525 1632 531
rect -108 519 -81 525
rect -75 519 15 525
rect 21 519 63 525
rect 69 519 111 525
rect 117 519 159 525
rect 165 519 207 525
rect 213 519 255 525
rect 261 519 303 525
rect 309 519 351 525
rect 357 519 399 525
rect 405 519 447 525
rect 453 519 495 525
rect 501 519 543 525
rect 549 519 591 525
rect 597 519 639 525
rect 645 519 687 525
rect 693 519 735 525
rect 741 519 783 525
rect 789 519 831 525
rect 837 519 879 525
rect 885 519 927 525
rect 933 519 975 525
rect 981 519 1023 525
rect 1029 519 1071 525
rect 1077 519 1119 525
rect 1125 519 1167 525
rect 1173 519 1215 525
rect 1221 519 1263 525
rect 1269 519 1311 525
rect 1317 519 1359 525
rect 1365 519 1407 525
rect 1413 519 1455 525
rect 1461 519 1503 525
rect 1509 519 1599 525
rect 1605 519 1632 525
rect -108 516 1632 519
rect -108 477 1632 480
rect -108 471 -57 477
rect -51 471 -9 477
rect -3 471 39 477
rect 45 471 87 477
rect 93 471 135 477
rect 141 471 183 477
rect 189 471 231 477
rect 237 471 279 477
rect 285 471 327 477
rect 333 471 375 477
rect 381 471 423 477
rect 429 471 471 477
rect 477 471 519 477
rect 525 471 567 477
rect 573 471 615 477
rect 621 471 663 477
rect 669 471 711 477
rect 717 471 759 477
rect 765 471 807 477
rect 813 471 855 477
rect 861 471 903 477
rect 909 471 951 477
rect 957 471 999 477
rect 1005 471 1047 477
rect 1053 471 1095 477
rect 1101 471 1143 477
rect 1149 471 1191 477
rect 1197 471 1239 477
rect 1245 471 1287 477
rect 1293 471 1335 477
rect 1341 471 1383 477
rect 1389 471 1431 477
rect 1437 471 1479 477
rect 1485 471 1527 477
rect 1533 471 1575 477
rect 1581 471 1632 477
rect -108 462 1632 471
rect -108 453 1632 456
rect -108 447 -81 453
rect -75 447 -33 453
rect -27 447 15 453
rect 21 447 63 453
rect 69 447 111 453
rect 117 447 159 453
rect 165 447 207 453
rect 213 447 255 453
rect 261 447 303 453
rect 309 447 351 453
rect 357 447 399 453
rect 405 447 447 453
rect 453 447 495 453
rect 501 447 543 453
rect 549 447 591 453
rect 597 447 639 453
rect 645 447 687 453
rect 693 447 735 453
rect 741 447 783 453
rect 789 447 831 453
rect 837 447 879 453
rect 885 447 927 453
rect 933 447 975 453
rect 981 447 1023 453
rect 1029 447 1071 453
rect 1077 447 1119 453
rect 1125 447 1167 453
rect 1173 447 1215 453
rect 1221 447 1263 453
rect 1269 447 1311 453
rect 1317 447 1359 453
rect 1365 447 1407 453
rect 1413 447 1455 453
rect 1461 447 1503 453
rect 1509 447 1551 453
rect 1557 447 1599 453
rect 1605 447 1632 453
rect -108 444 1632 447
rect -108 429 1632 438
rect -108 423 -57 429
rect -51 423 -9 429
rect -3 423 39 429
rect 45 423 87 429
rect 93 423 183 429
rect 189 423 279 429
rect 285 423 375 429
rect 381 423 471 429
rect 477 423 567 429
rect 573 423 615 429
rect 621 423 663 429
rect 669 423 759 429
rect 765 423 855 429
rect 861 423 903 429
rect 909 423 951 429
rect 957 423 1047 429
rect 1053 423 1143 429
rect 1149 423 1239 429
rect 1245 423 1335 429
rect 1341 423 1431 429
rect 1437 423 1479 429
rect 1485 423 1527 429
rect 1533 423 1575 429
rect 1581 423 1632 429
rect -108 417 1632 423
rect -108 411 -57 417
rect -51 411 -9 417
rect -3 411 87 417
rect 93 411 183 417
rect 189 411 375 417
rect 381 411 567 417
rect 573 411 663 417
rect 669 411 759 417
rect 765 411 855 417
rect 861 411 951 417
rect 957 411 1143 417
rect 1149 411 1335 417
rect 1341 411 1431 417
rect 1437 411 1527 417
rect 1533 411 1575 417
rect 1581 411 1632 417
rect -108 405 1632 411
rect -108 399 -57 405
rect -51 399 -9 405
rect -3 399 87 405
rect 93 399 183 405
rect 189 399 375 405
rect 381 399 567 405
rect 573 399 663 405
rect 669 399 759 405
rect 765 399 855 405
rect 861 399 951 405
rect 957 399 1143 405
rect 1149 399 1335 405
rect 1341 399 1431 405
rect 1437 399 1527 405
rect 1533 399 1575 405
rect 1581 399 1632 405
rect -108 396 1632 399
rect 12 381 24 384
rect 12 375 15 381
rect 21 375 24 381
rect 12 372 24 375
rect 60 381 72 384
rect 60 375 63 381
rect 69 375 72 381
rect 60 372 72 375
rect 108 381 120 384
rect 108 375 111 381
rect 117 375 120 381
rect 108 372 120 375
rect 156 381 168 384
rect 156 375 159 381
rect 165 375 168 381
rect 156 372 168 375
rect 204 381 216 384
rect 204 375 207 381
rect 213 375 216 381
rect 204 372 216 375
rect 252 381 264 384
rect 252 375 255 381
rect 261 375 264 381
rect 252 372 264 375
rect 300 381 312 384
rect 300 375 303 381
rect 309 375 312 381
rect 300 372 312 375
rect 348 381 360 384
rect 348 375 351 381
rect 357 375 360 381
rect 348 372 360 375
rect 396 381 408 384
rect 396 375 399 381
rect 405 375 408 381
rect 396 372 408 375
rect 444 381 456 384
rect 444 375 447 381
rect 453 375 456 381
rect 444 372 456 375
rect 492 381 504 384
rect 492 375 495 381
rect 501 375 504 381
rect 492 372 504 375
rect 540 381 552 384
rect 540 375 543 381
rect 549 375 552 381
rect 540 372 552 375
rect 588 381 600 384
rect 588 375 591 381
rect 597 375 600 381
rect 588 372 600 375
rect 636 381 648 384
rect 636 375 639 381
rect 645 375 648 381
rect 636 372 648 375
rect 684 381 696 384
rect 684 375 687 381
rect 693 375 696 381
rect 684 372 696 375
rect 732 381 744 384
rect 732 375 735 381
rect 741 375 744 381
rect 732 372 744 375
rect 780 381 792 384
rect 780 375 783 381
rect 789 375 792 381
rect 780 372 792 375
rect 828 381 840 384
rect 828 375 831 381
rect 837 375 840 381
rect 828 372 840 375
rect 876 381 888 384
rect 876 375 879 381
rect 885 375 888 381
rect 876 372 888 375
rect 924 381 936 384
rect 924 375 927 381
rect 933 375 936 381
rect 924 372 936 375
rect 972 381 984 384
rect 972 375 975 381
rect 981 375 984 381
rect 972 372 984 375
rect 1020 381 1032 384
rect 1020 375 1023 381
rect 1029 375 1032 381
rect 1020 372 1032 375
rect 1068 381 1080 384
rect 1068 375 1071 381
rect 1077 375 1080 381
rect 1068 372 1080 375
rect 1116 381 1128 384
rect 1116 375 1119 381
rect 1125 375 1128 381
rect 1116 372 1128 375
rect 1164 381 1176 384
rect 1164 375 1167 381
rect 1173 375 1176 381
rect 1164 372 1176 375
rect 1212 381 1224 384
rect 1212 375 1215 381
rect 1221 375 1224 381
rect 1212 372 1224 375
rect 1260 381 1272 384
rect 1260 375 1263 381
rect 1269 375 1272 381
rect 1260 372 1272 375
rect 1308 381 1320 384
rect 1308 375 1311 381
rect 1317 375 1320 381
rect 1308 372 1320 375
rect 1356 381 1368 384
rect 1356 375 1359 381
rect 1365 375 1368 381
rect 1356 372 1368 375
rect 1404 381 1416 384
rect 1404 375 1407 381
rect 1413 375 1416 381
rect 1404 372 1416 375
rect 1452 381 1464 384
rect 1452 375 1455 381
rect 1461 375 1464 381
rect 1452 372 1464 375
rect 1500 381 1512 384
rect 1500 375 1503 381
rect 1509 375 1512 381
rect 1500 372 1512 375
rect -108 333 1632 336
rect -108 327 -57 333
rect -51 327 -9 333
rect -3 327 183 333
rect 189 327 375 333
rect 381 327 567 333
rect 573 327 759 333
rect 765 327 951 333
rect 957 327 1143 333
rect 1149 327 1335 333
rect 1341 327 1527 333
rect 1533 327 1575 333
rect 1581 327 1632 333
rect -108 324 1632 327
rect -108 309 1632 312
rect -108 303 495 309
rect 501 303 543 309
rect 549 303 975 309
rect 981 303 1023 309
rect 1029 303 1632 309
rect -108 300 1632 303
rect -108 285 1632 288
rect -108 279 -57 285
rect -51 279 -9 285
rect -3 279 183 285
rect 189 279 375 285
rect 381 279 567 285
rect 573 279 759 285
rect 765 279 951 285
rect 957 279 1143 285
rect 1149 279 1335 285
rect 1341 279 1527 285
rect 1533 279 1575 285
rect 1581 279 1632 285
rect -108 276 1632 279
rect -108 261 1632 264
rect -108 255 303 261
rect 309 255 351 261
rect 357 255 399 261
rect 405 255 447 261
rect 453 255 471 261
rect 477 255 1047 261
rect 1053 255 1071 261
rect 1077 255 1119 261
rect 1125 255 1167 261
rect 1173 255 1215 261
rect 1221 255 1632 261
rect -108 252 1632 255
rect -108 237 1632 240
rect -108 231 -57 237
rect -51 231 -9 237
rect -3 231 183 237
rect 189 231 375 237
rect 381 231 567 237
rect 573 231 759 237
rect 765 231 951 237
rect 957 231 1143 237
rect 1149 231 1335 237
rect 1341 231 1527 237
rect 1533 231 1575 237
rect 1581 231 1632 237
rect -108 228 1632 231
rect -108 213 1632 216
rect -108 207 207 213
rect 213 207 255 213
rect 261 207 1263 213
rect 1269 207 1311 213
rect 1317 207 1632 213
rect -108 204 1632 207
rect -108 189 1632 192
rect -108 183 -57 189
rect -51 183 -9 189
rect -3 183 183 189
rect 189 183 375 189
rect 381 183 567 189
rect 573 183 759 189
rect 765 183 951 189
rect 957 183 1143 189
rect 1149 183 1335 189
rect 1341 183 1527 189
rect 1533 183 1575 189
rect 1581 183 1632 189
rect -108 180 1632 183
rect -108 165 1632 168
rect -108 159 -81 165
rect -75 159 39 165
rect 45 159 135 165
rect 141 159 615 165
rect 621 159 711 165
rect 717 159 807 165
rect 813 159 903 165
rect 909 159 1383 165
rect 1389 159 1479 165
rect 1485 159 1599 165
rect 1605 159 1632 165
rect -108 150 1632 159
rect -108 141 1632 144
rect -108 135 15 141
rect 21 135 63 141
rect 69 135 111 141
rect 117 135 159 141
rect 165 135 279 141
rect 285 135 591 141
rect 597 135 639 141
rect 645 135 687 141
rect 693 135 735 141
rect 741 135 783 141
rect 789 135 831 141
rect 837 135 879 141
rect 885 135 927 141
rect 933 135 1239 141
rect 1245 135 1359 141
rect 1365 135 1407 141
rect 1413 135 1455 141
rect 1461 135 1503 141
rect 1509 135 1632 141
rect -108 132 1632 135
rect -108 117 1632 126
rect -108 111 -81 117
rect -75 111 39 117
rect 45 111 135 117
rect 141 111 615 117
rect 621 111 711 117
rect 717 111 807 117
rect 813 111 903 117
rect 909 111 1383 117
rect 1389 111 1479 117
rect 1485 111 1599 117
rect 1605 111 1632 117
rect -108 108 1632 111
rect -108 93 1632 96
rect -108 87 -57 93
rect -51 87 -9 93
rect -3 87 183 93
rect 189 87 375 93
rect 381 87 567 93
rect 573 87 759 93
rect 765 87 951 93
rect 957 87 1143 93
rect 1149 87 1335 93
rect 1341 87 1527 93
rect 1533 87 1575 93
rect 1581 87 1632 93
rect -108 84 1632 87
rect 12 69 24 72
rect 12 63 15 69
rect 21 63 24 69
rect 12 60 24 63
rect 60 69 72 72
rect 60 63 63 69
rect 69 63 72 69
rect 60 60 72 63
rect 108 69 120 72
rect 108 63 111 69
rect 117 63 120 69
rect 108 60 120 63
rect 156 69 168 72
rect 156 63 159 69
rect 165 63 168 69
rect 156 60 168 63
rect 204 69 216 72
rect 204 63 207 69
rect 213 63 216 69
rect 204 60 216 63
rect 252 69 264 72
rect 252 63 255 69
rect 261 63 264 69
rect 252 60 264 63
rect 300 69 312 72
rect 300 63 303 69
rect 309 63 312 69
rect 300 60 312 63
rect 348 69 360 72
rect 348 63 351 69
rect 357 63 360 69
rect 348 60 360 63
rect 396 69 408 72
rect 396 63 399 69
rect 405 63 408 69
rect 396 60 408 63
rect 444 69 456 72
rect 444 63 447 69
rect 453 63 456 69
rect 444 60 456 63
rect 492 69 504 72
rect 492 63 495 69
rect 501 63 504 69
rect 492 60 504 63
rect 540 69 552 72
rect 540 63 543 69
rect 549 63 552 69
rect 540 60 552 63
rect 588 69 600 72
rect 588 63 591 69
rect 597 63 600 69
rect 588 60 600 63
rect 636 69 648 72
rect 636 63 639 69
rect 645 63 648 69
rect 636 60 648 63
rect 684 69 696 72
rect 684 63 687 69
rect 693 63 696 69
rect 684 60 696 63
rect 732 69 744 72
rect 732 63 735 69
rect 741 63 744 69
rect 732 60 744 63
rect 780 69 792 72
rect 780 63 783 69
rect 789 63 792 69
rect 780 60 792 63
rect 828 69 840 72
rect 828 63 831 69
rect 837 63 840 69
rect 828 60 840 63
rect 876 69 888 72
rect 876 63 879 69
rect 885 63 888 69
rect 876 60 888 63
rect 924 69 936 72
rect 924 63 927 69
rect 933 63 936 69
rect 924 60 936 63
rect 972 69 984 72
rect 972 63 975 69
rect 981 63 984 69
rect 972 60 984 63
rect 1020 69 1032 72
rect 1020 63 1023 69
rect 1029 63 1032 69
rect 1020 60 1032 63
rect 1068 69 1080 72
rect 1068 63 1071 69
rect 1077 63 1080 69
rect 1068 60 1080 63
rect 1116 69 1128 72
rect 1116 63 1119 69
rect 1125 63 1128 69
rect 1116 60 1128 63
rect 1164 69 1176 72
rect 1164 63 1167 69
rect 1173 63 1176 69
rect 1164 60 1176 63
rect 1212 69 1224 72
rect 1212 63 1215 69
rect 1221 63 1224 69
rect 1212 60 1224 63
rect 1260 69 1272 72
rect 1260 63 1263 69
rect 1269 63 1272 69
rect 1260 60 1272 63
rect 1308 69 1320 72
rect 1308 63 1311 69
rect 1317 63 1320 69
rect 1308 60 1320 63
rect 1356 69 1368 72
rect 1356 63 1359 69
rect 1365 63 1368 69
rect 1356 60 1368 63
rect 1404 69 1416 72
rect 1404 63 1407 69
rect 1413 63 1416 69
rect 1404 60 1416 63
rect 1452 69 1464 72
rect 1452 63 1455 69
rect 1461 63 1464 69
rect 1452 60 1464 63
rect 1500 69 1512 72
rect 1500 63 1503 69
rect 1509 63 1512 69
rect 1500 60 1512 63
rect -108 45 1632 48
rect -108 39 -57 45
rect -51 39 -9 45
rect -3 39 87 45
rect 93 39 183 45
rect 189 39 375 45
rect 381 39 567 45
rect 573 39 663 45
rect 669 39 759 45
rect 765 39 855 45
rect 861 39 951 45
rect 957 39 1143 45
rect 1149 39 1335 45
rect 1341 39 1431 45
rect 1437 39 1527 45
rect 1533 39 1575 45
rect 1581 39 1632 45
rect -108 33 1632 39
rect -108 27 -57 33
rect -51 27 -9 33
rect -3 27 87 33
rect 93 27 183 33
rect 189 27 375 33
rect 381 27 567 33
rect 573 27 663 33
rect 669 27 759 33
rect 765 27 855 33
rect 861 27 951 33
rect 957 27 1143 33
rect 1149 27 1335 33
rect 1341 27 1431 33
rect 1437 27 1527 33
rect 1533 27 1575 33
rect 1581 27 1632 33
rect -108 21 1632 27
rect -108 15 -57 21
rect -51 15 -9 21
rect -3 15 87 21
rect 93 15 183 21
rect 189 15 375 21
rect 381 15 567 21
rect 573 15 663 21
rect 669 15 759 21
rect 765 15 855 21
rect 861 15 951 21
rect 957 15 1143 21
rect 1149 15 1335 21
rect 1341 15 1431 21
rect 1437 15 1527 21
rect 1533 15 1575 21
rect 1581 15 1632 21
rect -108 12 1632 15
<< via3 >>
rect 15 375 21 381
rect 63 375 69 381
rect 111 375 117 381
rect 159 375 165 381
rect 207 375 213 381
rect 255 375 261 381
rect 303 375 309 381
rect 351 375 357 381
rect 399 375 405 381
rect 447 375 453 381
rect 495 375 501 381
rect 543 375 549 381
rect 591 375 597 381
rect 639 375 645 381
rect 687 375 693 381
rect 735 375 741 381
rect 783 375 789 381
rect 831 375 837 381
rect 879 375 885 381
rect 927 375 933 381
rect 975 375 981 381
rect 1023 375 1029 381
rect 1071 375 1077 381
rect 1119 375 1125 381
rect 1167 375 1173 381
rect 1215 375 1221 381
rect 1263 375 1269 381
rect 1311 375 1317 381
rect 1359 375 1365 381
rect 1407 375 1413 381
rect 1455 375 1461 381
rect 1503 375 1509 381
rect 495 303 501 309
rect 543 303 549 309
rect 975 303 981 309
rect 1023 303 1029 309
rect 303 255 309 261
rect 351 255 357 261
rect 399 255 405 261
rect 447 255 453 261
rect 1071 255 1077 261
rect 1119 255 1125 261
rect 1167 255 1173 261
rect 1215 255 1221 261
rect 207 207 213 213
rect 255 207 261 213
rect 1263 207 1269 213
rect 1311 207 1317 213
rect -81 159 -75 165
rect 1599 159 1605 165
rect 15 135 21 141
rect 63 135 69 141
rect 111 135 117 141
rect 159 135 165 141
rect 591 135 597 141
rect 639 135 645 141
rect 687 135 693 141
rect 735 135 741 141
rect 783 135 789 141
rect 831 135 837 141
rect 879 135 885 141
rect 927 135 933 141
rect 1359 135 1365 141
rect 1407 135 1413 141
rect 1455 135 1461 141
rect 1503 135 1509 141
rect -81 111 -75 117
rect 1599 111 1605 117
rect 15 63 21 69
rect 63 63 69 69
rect 111 63 117 69
rect 159 63 165 69
rect 207 63 213 69
rect 255 63 261 69
rect 303 63 309 69
rect 351 63 357 69
rect 399 63 405 69
rect 447 63 453 69
rect 495 63 501 69
rect 543 63 549 69
rect 591 63 597 69
rect 639 63 645 69
rect 687 63 693 69
rect 735 63 741 69
rect 783 63 789 69
rect 831 63 837 69
rect 879 63 885 69
rect 927 63 933 69
rect 975 63 981 69
rect 1023 63 1029 69
rect 1071 63 1077 69
rect 1119 63 1125 69
rect 1167 63 1173 69
rect 1215 63 1221 69
rect 1263 63 1269 69
rect 1311 63 1317 69
rect 1359 63 1365 69
rect 1407 63 1413 69
rect 1455 63 1461 69
rect 1503 63 1509 69
<< metal4 >>
rect 12 381 24 384
rect 12 375 15 381
rect 21 375 24 381
rect 12 372 24 375
rect 60 381 72 384
rect 60 375 63 381
rect 69 375 72 381
rect 60 372 72 375
rect 108 381 120 384
rect 108 375 111 381
rect 117 375 120 381
rect 108 372 120 375
rect 156 381 168 384
rect 156 375 159 381
rect 165 375 168 381
rect 156 372 168 375
rect 204 381 216 384
rect 204 375 207 381
rect 213 375 216 381
rect 204 372 216 375
rect 252 381 264 384
rect 252 375 255 381
rect 261 375 264 381
rect 252 372 264 375
rect 300 381 312 384
rect 300 375 303 381
rect 309 375 312 381
rect 300 372 312 375
rect 348 381 360 384
rect 348 375 351 381
rect 357 375 360 381
rect 348 372 360 375
rect 396 381 408 384
rect 396 375 399 381
rect 405 375 408 381
rect 396 372 408 375
rect 444 381 456 384
rect 444 375 447 381
rect 453 375 456 381
rect 444 372 456 375
rect 492 381 504 384
rect 492 375 495 381
rect 501 375 504 381
rect 492 372 504 375
rect 540 381 552 384
rect 540 375 543 381
rect 549 375 552 381
rect 540 372 552 375
rect 588 381 600 384
rect 588 375 591 381
rect 597 375 600 381
rect 588 372 600 375
rect 636 381 648 384
rect 636 375 639 381
rect 645 375 648 381
rect 636 372 648 375
rect 684 381 696 384
rect 684 375 687 381
rect 693 375 696 381
rect 684 372 696 375
rect 732 381 744 384
rect 732 375 735 381
rect 741 375 744 381
rect 732 372 744 375
rect 780 381 792 384
rect 780 375 783 381
rect 789 375 792 381
rect 780 372 792 375
rect 828 381 840 384
rect 828 375 831 381
rect 837 375 840 381
rect 828 372 840 375
rect 876 381 888 384
rect 876 375 879 381
rect 885 375 888 381
rect 876 372 888 375
rect 924 381 936 384
rect 924 375 927 381
rect 933 375 936 381
rect 924 372 936 375
rect 972 381 984 384
rect 972 375 975 381
rect 981 375 984 381
rect 972 372 984 375
rect 1020 381 1032 384
rect 1020 375 1023 381
rect 1029 375 1032 381
rect 1020 372 1032 375
rect 1068 381 1080 384
rect 1068 375 1071 381
rect 1077 375 1080 381
rect 1068 372 1080 375
rect 1116 381 1128 384
rect 1116 375 1119 381
rect 1125 375 1128 381
rect 1116 372 1128 375
rect 1164 381 1176 384
rect 1164 375 1167 381
rect 1173 375 1176 381
rect 1164 372 1176 375
rect 1212 381 1224 384
rect 1212 375 1215 381
rect 1221 375 1224 381
rect 1212 372 1224 375
rect 1260 381 1272 384
rect 1260 375 1263 381
rect 1269 375 1272 381
rect 1260 372 1272 375
rect 1308 381 1320 384
rect 1308 375 1311 381
rect 1317 375 1320 381
rect 1308 372 1320 375
rect 1356 381 1368 384
rect 1356 375 1359 381
rect 1365 375 1368 381
rect 1356 372 1368 375
rect 1404 381 1416 384
rect 1404 375 1407 381
rect 1413 375 1416 381
rect 1404 372 1416 375
rect 1452 381 1464 384
rect 1452 375 1455 381
rect 1461 375 1464 381
rect 1452 372 1464 375
rect 1500 381 1512 384
rect 1500 375 1503 381
rect 1509 375 1512 381
rect 1500 372 1512 375
rect 492 309 504 312
rect 492 303 495 309
rect 501 303 504 309
rect 492 300 504 303
rect 540 309 552 312
rect 540 303 543 309
rect 549 303 552 309
rect 540 300 552 303
rect 972 309 984 312
rect 972 303 975 309
rect 981 303 984 309
rect 972 300 984 303
rect 1020 309 1032 312
rect 1020 303 1023 309
rect 1029 303 1032 309
rect 1020 300 1032 303
rect 300 261 312 264
rect 300 255 303 261
rect 309 255 312 261
rect 300 252 312 255
rect 348 261 360 264
rect 348 255 351 261
rect 357 255 360 261
rect 348 252 360 255
rect 396 261 408 264
rect 396 255 399 261
rect 405 255 408 261
rect 396 252 408 255
rect 444 261 456 264
rect 444 255 447 261
rect 453 255 456 261
rect 444 252 456 255
rect 1068 261 1080 264
rect 1068 255 1071 261
rect 1077 255 1080 261
rect 1068 252 1080 255
rect 1116 261 1128 264
rect 1116 255 1119 261
rect 1125 255 1128 261
rect 1116 252 1128 255
rect 1164 261 1176 264
rect 1164 255 1167 261
rect 1173 255 1176 261
rect 1164 252 1176 255
rect 1212 261 1224 264
rect 1212 255 1215 261
rect 1221 255 1224 261
rect 1212 252 1224 255
rect 204 213 216 216
rect 204 207 207 213
rect 213 207 216 213
rect 204 204 216 207
rect 252 213 264 216
rect 252 207 255 213
rect 261 207 264 213
rect 252 204 264 207
rect 1260 213 1272 216
rect 1260 207 1263 213
rect 1269 207 1272 213
rect 1260 204 1272 207
rect 1308 213 1320 216
rect 1308 207 1311 213
rect 1317 207 1320 213
rect 1308 204 1320 207
rect -108 144 -96 168
rect -84 165 -72 168
rect -84 159 -81 165
rect -75 159 -72 165
rect -84 117 -72 159
rect 1596 165 1608 168
rect 1596 159 1599 165
rect 1605 159 1608 165
rect 12 141 24 144
rect 12 135 15 141
rect 21 135 24 141
rect 12 132 24 135
rect 60 141 72 144
rect 60 135 63 141
rect 69 135 72 141
rect 60 132 72 135
rect 108 141 120 144
rect 108 135 111 141
rect 117 135 120 141
rect 108 132 120 135
rect 156 141 168 144
rect 156 135 159 141
rect 165 135 168 141
rect 156 132 168 135
rect 588 141 600 144
rect 588 135 591 141
rect 597 135 600 141
rect 588 132 600 135
rect 636 141 648 144
rect 636 135 639 141
rect 645 135 648 141
rect 636 132 648 135
rect 684 141 696 144
rect 684 135 687 141
rect 693 135 696 141
rect 684 132 696 135
rect 732 141 744 144
rect 732 135 735 141
rect 741 135 744 141
rect 732 132 744 135
rect 780 141 792 144
rect 780 135 783 141
rect 789 135 792 141
rect 780 132 792 135
rect 828 141 840 144
rect 828 135 831 141
rect 837 135 840 141
rect 828 132 840 135
rect 876 141 888 144
rect 876 135 879 141
rect 885 135 888 141
rect 876 132 888 135
rect 924 141 936 144
rect 924 135 927 141
rect 933 135 936 141
rect 924 132 936 135
rect 1356 141 1368 144
rect 1356 135 1359 141
rect 1365 135 1368 141
rect 1356 132 1368 135
rect 1404 141 1416 144
rect 1404 135 1407 141
rect 1413 135 1416 141
rect 1404 132 1416 135
rect 1452 141 1464 144
rect 1452 135 1455 141
rect 1461 135 1464 141
rect 1452 132 1464 135
rect 1500 141 1512 144
rect 1500 135 1503 141
rect 1509 135 1512 141
rect 1500 132 1512 135
rect -84 111 -81 117
rect -75 111 -72 117
rect -84 -171 -72 111
rect 1596 117 1608 159
rect 1620 144 1632 168
rect 1596 111 1599 117
rect 1605 111 1608 117
rect 12 69 24 72
rect 12 63 15 69
rect 21 63 24 69
rect 12 60 24 63
rect 60 69 72 72
rect 60 63 63 69
rect 69 63 72 69
rect 60 60 72 63
rect 108 69 120 72
rect 108 63 111 69
rect 117 63 120 69
rect 108 60 120 63
rect 156 69 168 72
rect 156 63 159 69
rect 165 63 168 69
rect 156 60 168 63
rect 204 69 216 72
rect 204 63 207 69
rect 213 63 216 69
rect 204 60 216 63
rect 252 69 264 72
rect 252 63 255 69
rect 261 63 264 69
rect 252 60 264 63
rect 300 69 312 72
rect 300 63 303 69
rect 309 63 312 69
rect 300 60 312 63
rect 348 69 360 72
rect 348 63 351 69
rect 357 63 360 69
rect 348 60 360 63
rect 396 69 408 72
rect 396 63 399 69
rect 405 63 408 69
rect 396 60 408 63
rect 444 69 456 72
rect 444 63 447 69
rect 453 63 456 69
rect 444 60 456 63
rect 492 69 504 72
rect 492 63 495 69
rect 501 63 504 69
rect 492 60 504 63
rect 540 69 552 72
rect 540 63 543 69
rect 549 63 552 69
rect 540 60 552 63
rect 588 69 600 72
rect 588 63 591 69
rect 597 63 600 69
rect 588 60 600 63
rect 636 69 648 72
rect 636 63 639 69
rect 645 63 648 69
rect 636 60 648 63
rect 684 69 696 72
rect 684 63 687 69
rect 693 63 696 69
rect 684 60 696 63
rect 732 69 744 72
rect 732 63 735 69
rect 741 63 744 69
rect 732 60 744 63
rect 780 69 792 72
rect 780 63 783 69
rect 789 63 792 69
rect 780 60 792 63
rect 828 69 840 72
rect 828 63 831 69
rect 837 63 840 69
rect 828 60 840 63
rect 876 69 888 72
rect 876 63 879 69
rect 885 63 888 69
rect 876 60 888 63
rect 924 69 936 72
rect 924 63 927 69
rect 933 63 936 69
rect 924 60 936 63
rect 972 69 984 72
rect 972 63 975 69
rect 981 63 984 69
rect 972 60 984 63
rect 1020 69 1032 72
rect 1020 63 1023 69
rect 1029 63 1032 69
rect 1020 60 1032 63
rect 1068 69 1080 72
rect 1068 63 1071 69
rect 1077 63 1080 69
rect 1068 60 1080 63
rect 1116 69 1128 72
rect 1116 63 1119 69
rect 1125 63 1128 69
rect 1116 60 1128 63
rect 1164 69 1176 72
rect 1164 63 1167 69
rect 1173 63 1176 69
rect 1164 60 1176 63
rect 1212 69 1224 72
rect 1212 63 1215 69
rect 1221 63 1224 69
rect 1212 60 1224 63
rect 1260 69 1272 72
rect 1260 63 1263 69
rect 1269 63 1272 69
rect 1260 60 1272 63
rect 1308 69 1320 72
rect 1308 63 1311 69
rect 1317 63 1320 69
rect 1308 60 1320 63
rect 1356 69 1368 72
rect 1356 63 1359 69
rect 1365 63 1368 69
rect 1356 60 1368 63
rect 1404 69 1416 72
rect 1404 63 1407 69
rect 1413 63 1416 69
rect 1404 60 1416 63
rect 1452 69 1464 72
rect 1452 63 1455 69
rect 1461 63 1464 69
rect 1452 60 1464 63
rect 1500 69 1512 72
rect 1500 63 1503 69
rect 1509 63 1512 69
rect 1500 60 1512 63
rect -84 -177 -81 -171
rect -75 -177 -72 -171
rect -84 -180 -72 -177
rect -60 -27 1584 -24
rect -60 -33 -57 -27
rect -51 -33 -45 -27
rect -39 -33 -33 -27
rect -27 -33 -21 -27
rect -15 -33 -9 -27
rect -3 -33 3 -27
rect 9 -33 15 -27
rect 21 -33 27 -27
rect 33 -33 39 -27
rect 45 -33 51 -27
rect 57 -33 63 -27
rect 69 -33 75 -27
rect 81 -33 87 -27
rect 93 -33 99 -27
rect 105 -33 111 -27
rect 117 -33 123 -27
rect 129 -33 135 -27
rect 141 -33 147 -27
rect 153 -33 159 -27
rect 165 -33 171 -27
rect 177 -33 183 -27
rect 189 -33 195 -27
rect 201 -33 207 -27
rect 213 -33 219 -27
rect 225 -33 231 -27
rect 237 -33 243 -27
rect 249 -33 255 -27
rect 261 -33 267 -27
rect 273 -33 279 -27
rect 285 -33 291 -27
rect 297 -33 303 -27
rect 309 -33 315 -27
rect 321 -33 327 -27
rect 333 -33 339 -27
rect 345 -33 351 -27
rect 357 -33 363 -27
rect 369 -33 375 -27
rect 381 -33 387 -27
rect 393 -33 399 -27
rect 405 -33 411 -27
rect 417 -33 423 -27
rect 429 -33 435 -27
rect 441 -33 447 -27
rect 453 -33 459 -27
rect 465 -33 471 -27
rect 477 -33 483 -27
rect 489 -33 495 -27
rect 501 -33 507 -27
rect 513 -33 519 -27
rect 525 -33 531 -27
rect 537 -33 543 -27
rect 549 -33 555 -27
rect 561 -33 567 -27
rect 573 -33 579 -27
rect 585 -33 591 -27
rect 597 -33 603 -27
rect 609 -33 615 -27
rect 621 -33 627 -27
rect 633 -33 639 -27
rect 645 -33 651 -27
rect 657 -33 663 -27
rect 669 -33 675 -27
rect 681 -33 687 -27
rect 693 -33 699 -27
rect 705 -33 711 -27
rect 717 -33 723 -27
rect 729 -33 735 -27
rect 741 -33 747 -27
rect 753 -33 759 -27
rect 765 -33 771 -27
rect 777 -33 783 -27
rect 789 -33 795 -27
rect 801 -33 807 -27
rect 813 -33 819 -27
rect 825 -33 831 -27
rect 837 -33 843 -27
rect 849 -33 855 -27
rect 861 -33 867 -27
rect 873 -33 879 -27
rect 885 -33 891 -27
rect 897 -33 903 -27
rect 909 -33 915 -27
rect 921 -33 927 -27
rect 933 -33 939 -27
rect 945 -33 951 -27
rect 957 -33 963 -27
rect 969 -33 975 -27
rect 981 -33 987 -27
rect 993 -33 999 -27
rect 1005 -33 1011 -27
rect 1017 -33 1023 -27
rect 1029 -33 1035 -27
rect 1041 -33 1047 -27
rect 1053 -33 1059 -27
rect 1065 -33 1071 -27
rect 1077 -33 1083 -27
rect 1089 -33 1095 -27
rect 1101 -33 1107 -27
rect 1113 -33 1119 -27
rect 1125 -33 1131 -27
rect 1137 -33 1143 -27
rect 1149 -33 1155 -27
rect 1161 -33 1167 -27
rect 1173 -33 1179 -27
rect 1185 -33 1191 -27
rect 1197 -33 1203 -27
rect 1209 -33 1215 -27
rect 1221 -33 1227 -27
rect 1233 -33 1239 -27
rect 1245 -33 1251 -27
rect 1257 -33 1263 -27
rect 1269 -33 1275 -27
rect 1281 -33 1287 -27
rect 1293 -33 1299 -27
rect 1305 -33 1311 -27
rect 1317 -33 1323 -27
rect 1329 -33 1335 -27
rect 1341 -33 1347 -27
rect 1353 -33 1359 -27
rect 1365 -33 1371 -27
rect 1377 -33 1383 -27
rect 1389 -33 1395 -27
rect 1401 -33 1407 -27
rect 1413 -33 1419 -27
rect 1425 -33 1431 -27
rect 1437 -33 1443 -27
rect 1449 -33 1455 -27
rect 1461 -33 1467 -27
rect 1473 -33 1479 -27
rect 1485 -33 1491 -27
rect 1497 -33 1503 -27
rect 1509 -33 1515 -27
rect 1521 -33 1527 -27
rect 1533 -33 1539 -27
rect 1545 -33 1551 -27
rect 1557 -33 1563 -27
rect 1569 -33 1575 -27
rect 1581 -33 1584 -27
rect -60 -60 1584 -33
rect -60 -168 -48 -60
rect 1572 -168 1584 -60
rect -60 -180 1584 -168
rect 1596 -171 1608 111
rect 1596 -177 1599 -171
rect 1605 -177 1608 -171
rect 1596 -180 1608 -177
<< via4 >>
rect 15 375 21 381
rect 63 375 69 381
rect 111 375 117 381
rect 159 375 165 381
rect 207 375 213 381
rect 255 375 261 381
rect 303 375 309 381
rect 351 375 357 381
rect 399 375 405 381
rect 447 375 453 381
rect 495 375 501 381
rect 543 375 549 381
rect 591 375 597 381
rect 639 375 645 381
rect 687 375 693 381
rect 735 375 741 381
rect 783 375 789 381
rect 831 375 837 381
rect 879 375 885 381
rect 927 375 933 381
rect 975 375 981 381
rect 1023 375 1029 381
rect 1071 375 1077 381
rect 1119 375 1125 381
rect 1167 375 1173 381
rect 1215 375 1221 381
rect 1263 375 1269 381
rect 1311 375 1317 381
rect 1359 375 1365 381
rect 1407 375 1413 381
rect 1455 375 1461 381
rect 1503 375 1509 381
rect 495 303 501 309
rect 543 303 549 309
rect 975 303 981 309
rect 1023 303 1029 309
rect 303 255 309 261
rect 351 255 357 261
rect 399 255 405 261
rect 447 255 453 261
rect 1071 255 1077 261
rect 1119 255 1125 261
rect 1167 255 1173 261
rect 1215 255 1221 261
rect 207 207 213 213
rect 255 207 261 213
rect 1263 207 1269 213
rect 1311 207 1317 213
rect 15 135 21 141
rect 63 135 69 141
rect 111 135 117 141
rect 159 135 165 141
rect 591 135 597 141
rect 639 135 645 141
rect 687 135 693 141
rect 735 135 741 141
rect 783 135 789 141
rect 831 135 837 141
rect 879 135 885 141
rect 927 135 933 141
rect 1359 135 1365 141
rect 1407 135 1413 141
rect 1455 135 1461 141
rect 1503 135 1509 141
rect 15 63 21 69
rect 63 63 69 69
rect 111 63 117 69
rect 159 63 165 69
rect 207 63 213 69
rect 255 63 261 69
rect 303 63 309 69
rect 351 63 357 69
rect 399 63 405 69
rect 447 63 453 69
rect 495 63 501 69
rect 543 63 549 69
rect 591 63 597 69
rect 639 63 645 69
rect 687 63 693 69
rect 735 63 741 69
rect 783 63 789 69
rect 831 63 837 69
rect 879 63 885 69
rect 927 63 933 69
rect 975 63 981 69
rect 1023 63 1029 69
rect 1071 63 1077 69
rect 1119 63 1125 69
rect 1167 63 1173 69
rect 1215 63 1221 69
rect 1263 63 1269 69
rect 1311 63 1317 69
rect 1359 63 1365 69
rect 1407 63 1413 69
rect 1455 63 1461 69
rect 1503 63 1509 69
rect -81 -177 -75 -171
rect -57 -33 -51 -27
rect -45 -33 -39 -27
rect -33 -33 -27 -27
rect -21 -33 -15 -27
rect -9 -33 -3 -27
rect 3 -33 9 -27
rect 15 -33 21 -27
rect 27 -33 33 -27
rect 39 -33 45 -27
rect 51 -33 57 -27
rect 63 -33 69 -27
rect 75 -33 81 -27
rect 87 -33 93 -27
rect 99 -33 105 -27
rect 111 -33 117 -27
rect 123 -33 129 -27
rect 135 -33 141 -27
rect 147 -33 153 -27
rect 159 -33 165 -27
rect 171 -33 177 -27
rect 183 -33 189 -27
rect 195 -33 201 -27
rect 207 -33 213 -27
rect 219 -33 225 -27
rect 231 -33 237 -27
rect 243 -33 249 -27
rect 255 -33 261 -27
rect 267 -33 273 -27
rect 279 -33 285 -27
rect 291 -33 297 -27
rect 303 -33 309 -27
rect 315 -33 321 -27
rect 327 -33 333 -27
rect 339 -33 345 -27
rect 351 -33 357 -27
rect 363 -33 369 -27
rect 375 -33 381 -27
rect 387 -33 393 -27
rect 399 -33 405 -27
rect 411 -33 417 -27
rect 423 -33 429 -27
rect 435 -33 441 -27
rect 447 -33 453 -27
rect 459 -33 465 -27
rect 471 -33 477 -27
rect 483 -33 489 -27
rect 495 -33 501 -27
rect 507 -33 513 -27
rect 519 -33 525 -27
rect 531 -33 537 -27
rect 543 -33 549 -27
rect 555 -33 561 -27
rect 567 -33 573 -27
rect 579 -33 585 -27
rect 591 -33 597 -27
rect 603 -33 609 -27
rect 615 -33 621 -27
rect 627 -33 633 -27
rect 639 -33 645 -27
rect 651 -33 657 -27
rect 663 -33 669 -27
rect 675 -33 681 -27
rect 687 -33 693 -27
rect 699 -33 705 -27
rect 711 -33 717 -27
rect 723 -33 729 -27
rect 735 -33 741 -27
rect 747 -33 753 -27
rect 759 -33 765 -27
rect 771 -33 777 -27
rect 783 -33 789 -27
rect 795 -33 801 -27
rect 807 -33 813 -27
rect 819 -33 825 -27
rect 831 -33 837 -27
rect 843 -33 849 -27
rect 855 -33 861 -27
rect 867 -33 873 -27
rect 879 -33 885 -27
rect 891 -33 897 -27
rect 903 -33 909 -27
rect 915 -33 921 -27
rect 927 -33 933 -27
rect 939 -33 945 -27
rect 951 -33 957 -27
rect 963 -33 969 -27
rect 975 -33 981 -27
rect 987 -33 993 -27
rect 999 -33 1005 -27
rect 1011 -33 1017 -27
rect 1023 -33 1029 -27
rect 1035 -33 1041 -27
rect 1047 -33 1053 -27
rect 1059 -33 1065 -27
rect 1071 -33 1077 -27
rect 1083 -33 1089 -27
rect 1095 -33 1101 -27
rect 1107 -33 1113 -27
rect 1119 -33 1125 -27
rect 1131 -33 1137 -27
rect 1143 -33 1149 -27
rect 1155 -33 1161 -27
rect 1167 -33 1173 -27
rect 1179 -33 1185 -27
rect 1191 -33 1197 -27
rect 1203 -33 1209 -27
rect 1215 -33 1221 -27
rect 1227 -33 1233 -27
rect 1239 -33 1245 -27
rect 1251 -33 1257 -27
rect 1263 -33 1269 -27
rect 1275 -33 1281 -27
rect 1287 -33 1293 -27
rect 1299 -33 1305 -27
rect 1311 -33 1317 -27
rect 1323 -33 1329 -27
rect 1335 -33 1341 -27
rect 1347 -33 1353 -27
rect 1359 -33 1365 -27
rect 1371 -33 1377 -27
rect 1383 -33 1389 -27
rect 1395 -33 1401 -27
rect 1407 -33 1413 -27
rect 1419 -33 1425 -27
rect 1431 -33 1437 -27
rect 1443 -33 1449 -27
rect 1455 -33 1461 -27
rect 1467 -33 1473 -27
rect 1479 -33 1485 -27
rect 1491 -33 1497 -27
rect 1503 -33 1509 -27
rect 1515 -33 1521 -27
rect 1527 -33 1533 -27
rect 1539 -33 1545 -27
rect 1551 -33 1557 -27
rect 1563 -33 1569 -27
rect 1575 -33 1581 -27
rect 1599 -177 1605 -171
<< metal5 >>
rect 12 381 24 384
rect 12 375 15 381
rect 21 375 24 381
rect 12 141 24 375
rect 12 135 15 141
rect 21 135 24 141
rect 12 69 24 135
rect 12 63 15 69
rect 21 63 24 69
rect 12 60 24 63
rect 60 381 72 384
rect 60 375 63 381
rect 69 375 72 381
rect 60 141 72 375
rect 60 135 63 141
rect 69 135 72 141
rect 60 69 72 135
rect 60 63 63 69
rect 69 63 72 69
rect 60 -24 72 63
rect 108 381 120 384
rect 108 375 111 381
rect 117 375 120 381
rect 108 141 120 375
rect 108 135 111 141
rect 117 135 120 141
rect 108 69 120 135
rect 108 63 111 69
rect 117 63 120 69
rect 108 -24 120 63
rect 156 381 168 384
rect 156 375 159 381
rect 165 375 168 381
rect 156 141 168 375
rect 156 135 159 141
rect 165 135 168 141
rect 156 69 168 135
rect 156 63 159 69
rect 165 63 168 69
rect 156 60 168 63
rect 204 381 216 384
rect 204 375 207 381
rect 213 375 216 381
rect 204 213 216 375
rect 204 207 207 213
rect 213 207 216 213
rect 204 69 216 207
rect 204 63 207 69
rect 213 63 216 69
rect 204 60 216 63
rect 252 381 264 384
rect 252 375 255 381
rect 261 375 264 381
rect 252 213 264 375
rect 252 207 255 213
rect 261 207 264 213
rect 252 69 264 207
rect 252 63 255 69
rect 261 63 264 69
rect 252 60 264 63
rect 300 381 312 384
rect 300 375 303 381
rect 309 375 312 381
rect 300 261 312 375
rect 300 255 303 261
rect 309 255 312 261
rect 300 69 312 255
rect 300 63 303 69
rect 309 63 312 69
rect 300 60 312 63
rect 348 381 360 384
rect 348 375 351 381
rect 357 375 360 381
rect 348 261 360 375
rect 348 255 351 261
rect 357 255 360 261
rect 348 69 360 255
rect 348 63 351 69
rect 357 63 360 69
rect 348 60 360 63
rect 396 381 408 384
rect 396 375 399 381
rect 405 375 408 381
rect 396 261 408 375
rect 396 255 399 261
rect 405 255 408 261
rect 396 69 408 255
rect 396 63 399 69
rect 405 63 408 69
rect 396 60 408 63
rect 444 381 456 384
rect 444 375 447 381
rect 453 375 456 381
rect 444 261 456 375
rect 444 255 447 261
rect 453 255 456 261
rect 444 69 456 255
rect 444 63 447 69
rect 453 63 456 69
rect 444 60 456 63
rect 492 381 504 384
rect 492 375 495 381
rect 501 375 504 381
rect 492 309 504 375
rect 492 303 495 309
rect 501 303 504 309
rect 492 69 504 303
rect 492 63 495 69
rect 501 63 504 69
rect 492 60 504 63
rect 540 381 552 384
rect 540 375 543 381
rect 549 375 552 381
rect 540 309 552 375
rect 540 303 543 309
rect 549 303 552 309
rect 540 69 552 303
rect 540 63 543 69
rect 549 63 552 69
rect 540 60 552 63
rect 588 381 600 384
rect 588 375 591 381
rect 597 375 600 381
rect 588 141 600 375
rect 588 135 591 141
rect 597 135 600 141
rect 588 69 600 135
rect 588 63 591 69
rect 597 63 600 69
rect 588 60 600 63
rect 636 381 648 384
rect 636 375 639 381
rect 645 375 648 381
rect 636 141 648 375
rect 636 135 639 141
rect 645 135 648 141
rect 636 69 648 135
rect 636 63 639 69
rect 645 63 648 69
rect 636 -24 648 63
rect 684 381 696 384
rect 684 375 687 381
rect 693 375 696 381
rect 684 141 696 375
rect 684 135 687 141
rect 693 135 696 141
rect 684 69 696 135
rect 684 63 687 69
rect 693 63 696 69
rect 684 -24 696 63
rect 732 381 744 384
rect 732 375 735 381
rect 741 375 744 381
rect 732 141 744 375
rect 732 135 735 141
rect 741 135 744 141
rect 732 69 744 135
rect 732 63 735 69
rect 741 63 744 69
rect 732 60 744 63
rect 780 381 792 384
rect 780 375 783 381
rect 789 375 792 381
rect 780 141 792 375
rect 780 135 783 141
rect 789 135 792 141
rect 780 69 792 135
rect 780 63 783 69
rect 789 63 792 69
rect 780 60 792 63
rect 828 381 840 384
rect 828 375 831 381
rect 837 375 840 381
rect 828 141 840 375
rect 828 135 831 141
rect 837 135 840 141
rect 828 69 840 135
rect 828 63 831 69
rect 837 63 840 69
rect 828 -24 840 63
rect 876 381 888 384
rect 876 375 879 381
rect 885 375 888 381
rect 876 141 888 375
rect 876 135 879 141
rect 885 135 888 141
rect 876 69 888 135
rect 876 63 879 69
rect 885 63 888 69
rect 876 -24 888 63
rect 924 381 936 384
rect 924 375 927 381
rect 933 375 936 381
rect 924 141 936 375
rect 924 135 927 141
rect 933 135 936 141
rect 924 69 936 135
rect 924 63 927 69
rect 933 63 936 69
rect 924 60 936 63
rect 972 381 984 384
rect 972 375 975 381
rect 981 375 984 381
rect 972 309 984 375
rect 972 303 975 309
rect 981 303 984 309
rect 972 69 984 303
rect 972 63 975 69
rect 981 63 984 69
rect 972 60 984 63
rect 1020 381 1032 384
rect 1020 375 1023 381
rect 1029 375 1032 381
rect 1020 309 1032 375
rect 1020 303 1023 309
rect 1029 303 1032 309
rect 1020 69 1032 303
rect 1020 63 1023 69
rect 1029 63 1032 69
rect 1020 60 1032 63
rect 1068 381 1080 384
rect 1068 375 1071 381
rect 1077 375 1080 381
rect 1068 261 1080 375
rect 1068 255 1071 261
rect 1077 255 1080 261
rect 1068 69 1080 255
rect 1068 63 1071 69
rect 1077 63 1080 69
rect 1068 60 1080 63
rect 1116 381 1128 384
rect 1116 375 1119 381
rect 1125 375 1128 381
rect 1116 261 1128 375
rect 1116 255 1119 261
rect 1125 255 1128 261
rect 1116 69 1128 255
rect 1116 63 1119 69
rect 1125 63 1128 69
rect 1116 60 1128 63
rect 1164 381 1176 384
rect 1164 375 1167 381
rect 1173 375 1176 381
rect 1164 261 1176 375
rect 1164 255 1167 261
rect 1173 255 1176 261
rect 1164 69 1176 255
rect 1164 63 1167 69
rect 1173 63 1176 69
rect 1164 60 1176 63
rect 1212 381 1224 384
rect 1212 375 1215 381
rect 1221 375 1224 381
rect 1212 261 1224 375
rect 1212 255 1215 261
rect 1221 255 1224 261
rect 1212 69 1224 255
rect 1212 63 1215 69
rect 1221 63 1224 69
rect 1212 60 1224 63
rect 1260 381 1272 384
rect 1260 375 1263 381
rect 1269 375 1272 381
rect 1260 213 1272 375
rect 1260 207 1263 213
rect 1269 207 1272 213
rect 1260 69 1272 207
rect 1260 63 1263 69
rect 1269 63 1272 69
rect 1260 60 1272 63
rect 1308 381 1320 384
rect 1308 375 1311 381
rect 1317 375 1320 381
rect 1308 213 1320 375
rect 1308 207 1311 213
rect 1317 207 1320 213
rect 1308 69 1320 207
rect 1308 63 1311 69
rect 1317 63 1320 69
rect 1308 60 1320 63
rect 1356 381 1368 384
rect 1356 375 1359 381
rect 1365 375 1368 381
rect 1356 141 1368 375
rect 1356 135 1359 141
rect 1365 135 1368 141
rect 1356 69 1368 135
rect 1356 63 1359 69
rect 1365 63 1368 69
rect 1356 60 1368 63
rect 1404 381 1416 384
rect 1404 375 1407 381
rect 1413 375 1416 381
rect 1404 141 1416 375
rect 1404 135 1407 141
rect 1413 135 1416 141
rect 1404 69 1416 135
rect 1404 63 1407 69
rect 1413 63 1416 69
rect 1404 -24 1416 63
rect 1452 381 1464 384
rect 1452 375 1455 381
rect 1461 375 1464 381
rect 1452 141 1464 375
rect 1452 135 1455 141
rect 1461 135 1464 141
rect 1452 69 1464 135
rect 1452 63 1455 69
rect 1461 63 1464 69
rect 1452 -24 1464 63
rect 1500 381 1512 384
rect 1500 375 1503 381
rect 1509 375 1512 381
rect 1500 141 1512 375
rect 1500 135 1503 141
rect 1509 135 1512 141
rect 1500 69 1512 135
rect 1500 63 1503 69
rect 1509 63 1512 69
rect 1500 60 1512 63
rect -60 -27 1584 -24
rect -60 -33 -57 -27
rect -51 -33 -45 -27
rect -39 -33 -33 -27
rect -27 -33 -21 -27
rect -15 -33 -9 -27
rect -3 -33 3 -27
rect 9 -33 15 -27
rect 21 -33 27 -27
rect 33 -33 39 -27
rect 45 -33 51 -27
rect 57 -33 63 -27
rect 69 -33 75 -27
rect 81 -33 87 -27
rect 93 -33 99 -27
rect 105 -33 111 -27
rect 117 -33 123 -27
rect 129 -33 135 -27
rect 141 -33 147 -27
rect 153 -33 159 -27
rect 165 -33 171 -27
rect 177 -33 183 -27
rect 189 -33 195 -27
rect 201 -33 207 -27
rect 213 -33 219 -27
rect 225 -33 231 -27
rect 237 -33 243 -27
rect 249 -33 255 -27
rect 261 -33 267 -27
rect 273 -33 279 -27
rect 285 -33 291 -27
rect 297 -33 303 -27
rect 309 -33 315 -27
rect 321 -33 327 -27
rect 333 -33 339 -27
rect 345 -33 351 -27
rect 357 -33 363 -27
rect 369 -33 375 -27
rect 381 -33 387 -27
rect 393 -33 399 -27
rect 405 -33 411 -27
rect 417 -33 423 -27
rect 429 -33 435 -27
rect 441 -33 447 -27
rect 453 -33 459 -27
rect 465 -33 471 -27
rect 477 -33 483 -27
rect 489 -33 495 -27
rect 501 -33 507 -27
rect 513 -33 519 -27
rect 525 -33 531 -27
rect 537 -33 543 -27
rect 549 -33 555 -27
rect 561 -33 567 -27
rect 573 -33 579 -27
rect 585 -33 591 -27
rect 597 -33 603 -27
rect 609 -33 615 -27
rect 621 -33 627 -27
rect 633 -33 639 -27
rect 645 -33 651 -27
rect 657 -33 663 -27
rect 669 -33 675 -27
rect 681 -33 687 -27
rect 693 -33 699 -27
rect 705 -33 711 -27
rect 717 -33 723 -27
rect 729 -33 735 -27
rect 741 -33 747 -27
rect 753 -33 759 -27
rect 765 -33 771 -27
rect 777 -33 783 -27
rect 789 -33 795 -27
rect 801 -33 807 -27
rect 813 -33 819 -27
rect 825 -33 831 -27
rect 837 -33 843 -27
rect 849 -33 855 -27
rect 861 -33 867 -27
rect 873 -33 879 -27
rect 885 -33 891 -27
rect 897 -33 903 -27
rect 909 -33 915 -27
rect 921 -33 927 -27
rect 933 -33 939 -27
rect 945 -33 951 -27
rect 957 -33 963 -27
rect 969 -33 975 -27
rect 981 -33 987 -27
rect 993 -33 999 -27
rect 1005 -33 1011 -27
rect 1017 -33 1023 -27
rect 1029 -33 1035 -27
rect 1041 -33 1047 -27
rect 1053 -33 1059 -27
rect 1065 -33 1071 -27
rect 1077 -33 1083 -27
rect 1089 -33 1095 -27
rect 1101 -33 1107 -27
rect 1113 -33 1119 -27
rect 1125 -33 1131 -27
rect 1137 -33 1143 -27
rect 1149 -33 1155 -27
rect 1161 -33 1167 -27
rect 1173 -33 1179 -27
rect 1185 -33 1191 -27
rect 1197 -33 1203 -27
rect 1209 -33 1215 -27
rect 1221 -33 1227 -27
rect 1233 -33 1239 -27
rect 1245 -33 1251 -27
rect 1257 -33 1263 -27
rect 1269 -33 1275 -27
rect 1281 -33 1287 -27
rect 1293 -33 1299 -27
rect 1305 -33 1311 -27
rect 1317 -33 1323 -27
rect 1329 -33 1335 -27
rect 1341 -33 1347 -27
rect 1353 -33 1359 -27
rect 1365 -33 1371 -27
rect 1377 -33 1383 -27
rect 1389 -33 1395 -27
rect 1401 -33 1407 -27
rect 1413 -33 1419 -27
rect 1425 -33 1431 -27
rect 1437 -33 1443 -27
rect 1449 -33 1455 -27
rect 1461 -33 1467 -27
rect 1473 -33 1479 -27
rect 1485 -33 1491 -27
rect 1497 -33 1503 -27
rect 1509 -33 1515 -27
rect 1521 -33 1527 -27
rect 1533 -33 1539 -27
rect 1545 -33 1551 -27
rect 1557 -33 1563 -27
rect 1569 -33 1575 -27
rect 1581 -33 1584 -27
rect -60 -36 1584 -33
rect -60 -72 1584 -48
rect -60 -156 -36 -72
rect 1560 -156 1584 -72
rect -60 -168 1584 -156
rect -84 -171 1608 -168
rect -84 -177 -81 -171
rect -75 -177 1599 -171
rect 1605 -177 1608 -171
rect -84 -180 1608 -177
<< labels >>
rlabel metal3 -108 300 1632 312 0 im
port 1 nsew
rlabel metal3 -108 204 1632 216 0 ip
port 2 nsew
rlabel metal3 -108 156 1632 168 0 o
port 3 nsew
rlabel metal3 -108 588 1632 600 0 vdd
port 4 nsew
rlabel metal3 -108 564 1632 576 0 gp
port 5 nsew
rlabel metal3 -108 468 1632 480 0 vreg
port 6 nsew
rlabel metal3 -108 444 1632 456 0 bp
port 7 nsew
rlabel metal3 -108 24 1632 36 0 vss
port 8 nsew
rlabel metal3 -108 252 1632 264 0 x
rlabel metal3 -108 132 1632 144 0 y
<< end >>
