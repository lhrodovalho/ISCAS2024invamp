magic
tech gf180mcuC
timestamp 1697192518
<< nwell >>
rect -378 486 270 606
rect -378 342 270 462
<< nmos >>
rect -336 12 -324 48
rect -312 12 -300 48
rect -288 12 -276 48
rect -264 12 -252 48
rect -240 12 -228 48
rect -216 12 -204 48
rect -192 12 -180 48
rect -168 12 -156 48
rect -144 12 -132 48
rect -120 12 -108 48
rect -96 12 -84 48
rect -72 12 -60 48
rect -48 12 -36 48
rect -24 12 -12 48
rect 0 12 12 48
rect 24 12 36 48
rect 48 12 60 48
rect 72 12 84 48
rect 96 12 108 48
rect 120 12 132 48
rect 144 12 156 48
rect 168 12 180 48
rect 192 12 204 48
rect 216 12 228 48
<< pmos >>
rect -336 396 -324 426
rect -312 396 -300 426
rect -288 396 -276 426
rect -264 396 -252 426
rect -240 396 -228 426
rect -216 396 -204 426
rect -192 396 -180 426
rect -168 396 -156 426
rect -144 396 -132 426
rect -120 396 -108 426
rect -96 396 -84 426
rect -72 396 -60 426
rect -48 396 -36 426
rect -24 396 -12 426
rect 0 396 12 426
rect 24 396 36 426
rect 48 396 60 426
rect 72 396 84 426
rect 96 396 108 426
rect 120 396 132 426
rect 144 396 156 426
rect 168 396 180 426
rect 192 396 204 426
rect 216 396 228 426
<< mvpmos >>
rect -336 516 -324 552
rect -312 516 -300 552
rect -288 516 -276 552
rect -264 516 -252 552
rect -240 516 -228 552
rect -216 516 -204 552
rect -192 516 -180 552
rect -168 516 -156 552
rect -144 516 -132 552
rect -120 516 -108 552
rect -96 516 -84 552
rect -72 516 -60 552
rect -48 516 -36 552
rect -24 516 -12 552
rect 0 516 12 552
rect 24 516 36 552
rect 48 516 60 552
rect 72 516 84 552
rect 96 516 108 552
rect 120 516 132 552
rect 144 516 156 552
rect 168 516 180 552
rect 192 516 204 552
rect 216 516 228 552
<< ndiff >>
rect -348 45 -336 48
rect -348 39 -345 45
rect -339 39 -336 45
rect -348 33 -336 39
rect -348 27 -345 33
rect -339 27 -336 33
rect -348 21 -336 27
rect -348 15 -345 21
rect -339 15 -336 21
rect -348 12 -336 15
rect -324 45 -312 48
rect -324 39 -321 45
rect -315 39 -312 45
rect -324 33 -312 39
rect -324 27 -321 33
rect -315 27 -312 33
rect -324 21 -312 27
rect -324 15 -321 21
rect -315 15 -312 21
rect -324 12 -312 15
rect -300 45 -288 48
rect -300 39 -297 45
rect -291 39 -288 45
rect -300 33 -288 39
rect -300 27 -297 33
rect -291 27 -288 33
rect -300 21 -288 27
rect -300 15 -297 21
rect -291 15 -288 21
rect -300 12 -288 15
rect -276 45 -264 48
rect -276 39 -273 45
rect -267 39 -264 45
rect -276 33 -264 39
rect -276 27 -273 33
rect -267 27 -264 33
rect -276 21 -264 27
rect -276 15 -273 21
rect -267 15 -264 21
rect -276 12 -264 15
rect -252 45 -240 48
rect -252 39 -249 45
rect -243 39 -240 45
rect -252 33 -240 39
rect -252 27 -249 33
rect -243 27 -240 33
rect -252 21 -240 27
rect -252 15 -249 21
rect -243 15 -240 21
rect -252 12 -240 15
rect -228 45 -216 48
rect -228 39 -225 45
rect -219 39 -216 45
rect -228 33 -216 39
rect -228 27 -225 33
rect -219 27 -216 33
rect -228 21 -216 27
rect -228 15 -225 21
rect -219 15 -216 21
rect -228 12 -216 15
rect -204 45 -192 48
rect -204 39 -201 45
rect -195 39 -192 45
rect -204 33 -192 39
rect -204 27 -201 33
rect -195 27 -192 33
rect -204 21 -192 27
rect -204 15 -201 21
rect -195 15 -192 21
rect -204 12 -192 15
rect -180 45 -168 48
rect -180 39 -177 45
rect -171 39 -168 45
rect -180 33 -168 39
rect -180 27 -177 33
rect -171 27 -168 33
rect -180 21 -168 27
rect -180 15 -177 21
rect -171 15 -168 21
rect -180 12 -168 15
rect -156 45 -144 48
rect -156 39 -153 45
rect -147 39 -144 45
rect -156 33 -144 39
rect -156 27 -153 33
rect -147 27 -144 33
rect -156 21 -144 27
rect -156 15 -153 21
rect -147 15 -144 21
rect -156 12 -144 15
rect -132 45 -120 48
rect -132 39 -129 45
rect -123 39 -120 45
rect -132 33 -120 39
rect -132 27 -129 33
rect -123 27 -120 33
rect -132 21 -120 27
rect -132 15 -129 21
rect -123 15 -120 21
rect -132 12 -120 15
rect -108 45 -96 48
rect -108 39 -105 45
rect -99 39 -96 45
rect -108 33 -96 39
rect -108 27 -105 33
rect -99 27 -96 33
rect -108 21 -96 27
rect -108 15 -105 21
rect -99 15 -96 21
rect -108 12 -96 15
rect -84 12 -72 48
rect -60 45 -48 48
rect -60 39 -57 45
rect -51 39 -48 45
rect -60 33 -48 39
rect -60 27 -57 33
rect -51 27 -48 33
rect -60 21 -48 27
rect -60 15 -57 21
rect -51 15 -48 21
rect -60 12 -48 15
rect -36 12 -24 48
rect -12 45 0 48
rect -12 39 -9 45
rect -3 39 0 45
rect -12 33 0 39
rect -12 27 -9 33
rect -3 27 0 33
rect -12 21 0 27
rect -12 15 -9 21
rect -3 15 0 21
rect -12 12 0 15
rect 12 12 24 48
rect 36 45 48 48
rect 36 39 39 45
rect 45 39 48 45
rect 36 33 48 39
rect 36 27 39 33
rect 45 27 48 33
rect 36 21 48 27
rect 36 15 39 21
rect 45 15 48 21
rect 36 12 48 15
rect 60 12 72 48
rect 84 45 96 48
rect 84 39 87 45
rect 93 39 96 45
rect 84 33 96 39
rect 84 27 87 33
rect 93 27 96 33
rect 84 21 96 27
rect 84 15 87 21
rect 93 15 96 21
rect 84 12 96 15
rect 108 12 120 48
rect 132 45 144 48
rect 132 39 135 45
rect 141 39 144 45
rect 132 33 144 39
rect 132 27 135 33
rect 141 27 144 33
rect 132 21 144 27
rect 132 15 135 21
rect 141 15 144 21
rect 132 12 144 15
rect 156 12 168 48
rect 180 45 192 48
rect 180 39 183 45
rect 189 39 192 45
rect 180 33 192 39
rect 180 27 183 33
rect 189 27 192 33
rect 180 21 192 27
rect 180 15 183 21
rect 189 15 192 21
rect 180 12 192 15
rect 204 45 216 48
rect 204 39 207 45
rect 213 39 216 45
rect 204 33 216 39
rect 204 27 207 33
rect 213 27 216 33
rect 204 21 216 27
rect 204 15 207 21
rect 213 15 216 21
rect 204 12 216 15
rect 228 45 240 48
rect 228 39 231 45
rect 237 39 240 45
rect 228 33 240 39
rect 228 27 231 33
rect 237 27 240 33
rect 228 21 240 27
rect 228 15 231 21
rect 237 15 240 21
rect 228 12 240 15
<< pdiff >>
rect -348 417 -336 426
rect -348 411 -345 417
rect -339 411 -336 417
rect -348 405 -336 411
rect -348 399 -345 405
rect -339 399 -336 405
rect -348 396 -336 399
rect -324 417 -312 426
rect -324 411 -321 417
rect -315 411 -312 417
rect -324 405 -312 411
rect -324 399 -321 405
rect -315 399 -312 405
rect -324 396 -312 399
rect -300 417 -288 426
rect -300 411 -297 417
rect -291 411 -288 417
rect -300 405 -288 411
rect -300 399 -297 405
rect -291 399 -288 405
rect -300 396 -288 399
rect -276 417 -264 426
rect -276 411 -273 417
rect -267 411 -264 417
rect -276 405 -264 411
rect -276 399 -273 405
rect -267 399 -264 405
rect -276 396 -264 399
rect -252 417 -240 426
rect -252 411 -249 417
rect -243 411 -240 417
rect -252 405 -240 411
rect -252 399 -249 405
rect -243 399 -240 405
rect -252 396 -240 399
rect -228 417 -216 426
rect -228 411 -225 417
rect -219 411 -216 417
rect -228 405 -216 411
rect -228 399 -225 405
rect -219 399 -216 405
rect -228 396 -216 399
rect -204 417 -192 426
rect -204 411 -201 417
rect -195 411 -192 417
rect -204 405 -192 411
rect -204 399 -201 405
rect -195 399 -192 405
rect -204 396 -192 399
rect -180 417 -168 426
rect -180 411 -177 417
rect -171 411 -168 417
rect -180 405 -168 411
rect -180 399 -177 405
rect -171 399 -168 405
rect -180 396 -168 399
rect -156 417 -144 426
rect -156 411 -153 417
rect -147 411 -144 417
rect -156 405 -144 411
rect -156 399 -153 405
rect -147 399 -144 405
rect -156 396 -144 399
rect -132 417 -120 426
rect -132 411 -129 417
rect -123 411 -120 417
rect -132 405 -120 411
rect -132 399 -129 405
rect -123 399 -120 405
rect -132 396 -120 399
rect -108 417 -96 426
rect -108 411 -105 417
rect -99 411 -96 417
rect -108 405 -96 411
rect -108 399 -105 405
rect -99 399 -96 405
rect -108 396 -96 399
rect -84 417 -72 426
rect -84 411 -81 417
rect -75 411 -72 417
rect -84 405 -72 411
rect -84 399 -81 405
rect -75 399 -72 405
rect -84 396 -72 399
rect -60 417 -48 426
rect -60 411 -57 417
rect -51 411 -48 417
rect -60 405 -48 411
rect -60 399 -57 405
rect -51 399 -48 405
rect -60 396 -48 399
rect -36 417 -24 426
rect -36 411 -33 417
rect -27 411 -24 417
rect -36 405 -24 411
rect -36 399 -33 405
rect -27 399 -24 405
rect -36 396 -24 399
rect -12 417 0 426
rect -12 411 -9 417
rect -3 411 0 417
rect -12 405 0 411
rect -12 399 -9 405
rect -3 399 0 405
rect -12 396 0 399
rect 12 417 24 426
rect 12 411 15 417
rect 21 411 24 417
rect 12 405 24 411
rect 12 399 15 405
rect 21 399 24 405
rect 12 396 24 399
rect 36 417 48 426
rect 36 411 39 417
rect 45 411 48 417
rect 36 405 48 411
rect 36 399 39 405
rect 45 399 48 405
rect 36 396 48 399
rect 60 417 72 426
rect 60 411 63 417
rect 69 411 72 417
rect 60 405 72 411
rect 60 399 63 405
rect 69 399 72 405
rect 60 396 72 399
rect 84 417 96 426
rect 84 411 87 417
rect 93 411 96 417
rect 84 405 96 411
rect 84 399 87 405
rect 93 399 96 405
rect 84 396 96 399
rect 108 417 120 426
rect 108 411 111 417
rect 117 411 120 417
rect 108 405 120 411
rect 108 399 111 405
rect 117 399 120 405
rect 108 396 120 399
rect 132 417 144 426
rect 132 411 135 417
rect 141 411 144 417
rect 132 405 144 411
rect 132 399 135 405
rect 141 399 144 405
rect 132 396 144 399
rect 156 417 168 426
rect 156 411 159 417
rect 165 411 168 417
rect 156 405 168 411
rect 156 399 159 405
rect 165 399 168 405
rect 156 396 168 399
rect 180 417 192 426
rect 180 411 183 417
rect 189 411 192 417
rect 180 405 192 411
rect 180 399 183 405
rect 189 399 192 405
rect 180 396 192 399
rect 204 417 216 426
rect 204 411 207 417
rect 213 411 216 417
rect 204 405 216 411
rect 204 399 207 405
rect 213 399 216 405
rect 204 396 216 399
rect 228 417 240 426
rect 228 411 231 417
rect 237 411 240 417
rect 228 405 240 411
rect 228 399 231 405
rect 237 399 240 405
rect 228 396 240 399
<< mvpdiff >>
rect -348 549 -336 552
rect -348 543 -345 549
rect -339 543 -336 549
rect -348 537 -336 543
rect -348 531 -345 537
rect -339 531 -336 537
rect -348 525 -336 531
rect -348 519 -345 525
rect -339 519 -336 525
rect -348 516 -336 519
rect -324 549 -312 552
rect -324 543 -321 549
rect -315 543 -312 549
rect -324 537 -312 543
rect -324 531 -321 537
rect -315 531 -312 537
rect -324 525 -312 531
rect -324 519 -321 525
rect -315 519 -312 525
rect -324 516 -312 519
rect -300 549 -288 552
rect -300 543 -297 549
rect -291 543 -288 549
rect -300 537 -288 543
rect -300 531 -297 537
rect -291 531 -288 537
rect -300 525 -288 531
rect -300 519 -297 525
rect -291 519 -288 525
rect -300 516 -288 519
rect -276 549 -264 552
rect -276 543 -273 549
rect -267 543 -264 549
rect -276 537 -264 543
rect -276 531 -273 537
rect -267 531 -264 537
rect -276 525 -264 531
rect -276 519 -273 525
rect -267 519 -264 525
rect -276 516 -264 519
rect -252 549 -240 552
rect -252 543 -249 549
rect -243 543 -240 549
rect -252 537 -240 543
rect -252 531 -249 537
rect -243 531 -240 537
rect -252 525 -240 531
rect -252 519 -249 525
rect -243 519 -240 525
rect -252 516 -240 519
rect -228 549 -216 552
rect -228 543 -225 549
rect -219 543 -216 549
rect -228 537 -216 543
rect -228 531 -225 537
rect -219 531 -216 537
rect -228 525 -216 531
rect -228 519 -225 525
rect -219 519 -216 525
rect -228 516 -216 519
rect -204 549 -192 552
rect -204 543 -201 549
rect -195 543 -192 549
rect -204 537 -192 543
rect -204 531 -201 537
rect -195 531 -192 537
rect -204 525 -192 531
rect -204 519 -201 525
rect -195 519 -192 525
rect -204 516 -192 519
rect -180 549 -168 552
rect -180 543 -177 549
rect -171 543 -168 549
rect -180 537 -168 543
rect -180 531 -177 537
rect -171 531 -168 537
rect -180 525 -168 531
rect -180 519 -177 525
rect -171 519 -168 525
rect -180 516 -168 519
rect -156 549 -144 552
rect -156 543 -153 549
rect -147 543 -144 549
rect -156 537 -144 543
rect -156 531 -153 537
rect -147 531 -144 537
rect -156 525 -144 531
rect -156 519 -153 525
rect -147 519 -144 525
rect -156 516 -144 519
rect -132 549 -120 552
rect -132 543 -129 549
rect -123 543 -120 549
rect -132 537 -120 543
rect -132 531 -129 537
rect -123 531 -120 537
rect -132 525 -120 531
rect -132 519 -129 525
rect -123 519 -120 525
rect -132 516 -120 519
rect -108 549 -96 552
rect -108 543 -105 549
rect -99 543 -96 549
rect -108 537 -96 543
rect -108 531 -105 537
rect -99 531 -96 537
rect -108 525 -96 531
rect -108 519 -105 525
rect -99 519 -96 525
rect -108 516 -96 519
rect -84 549 -72 552
rect -84 543 -81 549
rect -75 543 -72 549
rect -84 537 -72 543
rect -84 531 -81 537
rect -75 531 -72 537
rect -84 525 -72 531
rect -84 519 -81 525
rect -75 519 -72 525
rect -84 516 -72 519
rect -60 549 -48 552
rect -60 543 -57 549
rect -51 543 -48 549
rect -60 537 -48 543
rect -60 531 -57 537
rect -51 531 -48 537
rect -60 525 -48 531
rect -60 519 -57 525
rect -51 519 -48 525
rect -60 516 -48 519
rect -36 549 -24 552
rect -36 543 -33 549
rect -27 543 -24 549
rect -36 537 -24 543
rect -36 531 -33 537
rect -27 531 -24 537
rect -36 525 -24 531
rect -36 519 -33 525
rect -27 519 -24 525
rect -36 516 -24 519
rect -12 549 0 552
rect -12 543 -9 549
rect -3 543 0 549
rect -12 537 0 543
rect -12 531 -9 537
rect -3 531 0 537
rect -12 525 0 531
rect -12 519 -9 525
rect -3 519 0 525
rect -12 516 0 519
rect 12 549 24 552
rect 12 543 15 549
rect 21 543 24 549
rect 12 537 24 543
rect 12 531 15 537
rect 21 531 24 537
rect 12 525 24 531
rect 12 519 15 525
rect 21 519 24 525
rect 12 516 24 519
rect 36 549 48 552
rect 36 543 39 549
rect 45 543 48 549
rect 36 537 48 543
rect 36 531 39 537
rect 45 531 48 537
rect 36 525 48 531
rect 36 519 39 525
rect 45 519 48 525
rect 36 516 48 519
rect 60 549 72 552
rect 60 543 63 549
rect 69 543 72 549
rect 60 537 72 543
rect 60 531 63 537
rect 69 531 72 537
rect 60 525 72 531
rect 60 519 63 525
rect 69 519 72 525
rect 60 516 72 519
rect 84 549 96 552
rect 84 543 87 549
rect 93 543 96 549
rect 84 537 96 543
rect 84 531 87 537
rect 93 531 96 537
rect 84 525 96 531
rect 84 519 87 525
rect 93 519 96 525
rect 84 516 96 519
rect 108 549 120 552
rect 108 543 111 549
rect 117 543 120 549
rect 108 537 120 543
rect 108 531 111 537
rect 117 531 120 537
rect 108 525 120 531
rect 108 519 111 525
rect 117 519 120 525
rect 108 516 120 519
rect 132 549 144 552
rect 132 543 135 549
rect 141 543 144 549
rect 132 537 144 543
rect 132 531 135 537
rect 141 531 144 537
rect 132 525 144 531
rect 132 519 135 525
rect 141 519 144 525
rect 132 516 144 519
rect 156 549 168 552
rect 156 543 159 549
rect 165 543 168 549
rect 156 537 168 543
rect 156 531 159 537
rect 165 531 168 537
rect 156 525 168 531
rect 156 519 159 525
rect 165 519 168 525
rect 156 516 168 519
rect 180 549 192 552
rect 180 543 183 549
rect 189 543 192 549
rect 180 537 192 543
rect 180 531 183 537
rect 189 531 192 537
rect 180 525 192 531
rect 180 519 183 525
rect 189 519 192 525
rect 180 516 192 519
rect 204 549 216 552
rect 204 543 207 549
rect 213 543 216 549
rect 204 537 216 543
rect 204 531 207 537
rect 213 531 216 537
rect 204 525 216 531
rect 204 519 207 525
rect 213 519 216 525
rect 204 516 216 519
rect 228 549 240 552
rect 228 543 231 549
rect 237 543 240 549
rect 228 537 240 543
rect 228 531 231 537
rect 237 531 240 537
rect 228 525 240 531
rect 228 519 231 525
rect 237 519 240 525
rect 228 516 240 519
<< ndiffc >>
rect -345 39 -339 45
rect -345 27 -339 33
rect -345 15 -339 21
rect -321 39 -315 45
rect -321 27 -315 33
rect -321 15 -315 21
rect -297 39 -291 45
rect -297 27 -291 33
rect -297 15 -291 21
rect -273 39 -267 45
rect -273 27 -267 33
rect -273 15 -267 21
rect -249 39 -243 45
rect -249 27 -243 33
rect -249 15 -243 21
rect -225 39 -219 45
rect -225 27 -219 33
rect -225 15 -219 21
rect -201 39 -195 45
rect -201 27 -195 33
rect -201 15 -195 21
rect -177 39 -171 45
rect -177 27 -171 33
rect -177 15 -171 21
rect -153 39 -147 45
rect -153 27 -147 33
rect -153 15 -147 21
rect -129 39 -123 45
rect -129 27 -123 33
rect -129 15 -123 21
rect -105 39 -99 45
rect -105 27 -99 33
rect -105 15 -99 21
rect -57 39 -51 45
rect -57 27 -51 33
rect -57 15 -51 21
rect -9 39 -3 45
rect -9 27 -3 33
rect -9 15 -3 21
rect 39 39 45 45
rect 39 27 45 33
rect 39 15 45 21
rect 87 39 93 45
rect 87 27 93 33
rect 87 15 93 21
rect 135 39 141 45
rect 135 27 141 33
rect 135 15 141 21
rect 183 39 189 45
rect 183 27 189 33
rect 183 15 189 21
rect 207 39 213 45
rect 207 27 213 33
rect 207 15 213 21
rect 231 39 237 45
rect 231 27 237 33
rect 231 15 237 21
<< pdiffc >>
rect -345 411 -339 417
rect -345 399 -339 405
rect -321 411 -315 417
rect -321 399 -315 405
rect -297 411 -291 417
rect -297 399 -291 405
rect -273 411 -267 417
rect -273 399 -267 405
rect -249 411 -243 417
rect -249 399 -243 405
rect -225 411 -219 417
rect -225 399 -219 405
rect -201 411 -195 417
rect -201 399 -195 405
rect -177 411 -171 417
rect -177 399 -171 405
rect -153 411 -147 417
rect -153 399 -147 405
rect -129 411 -123 417
rect -129 399 -123 405
rect -105 411 -99 417
rect -105 399 -99 405
rect -81 411 -75 417
rect -81 399 -75 405
rect -57 411 -51 417
rect -57 399 -51 405
rect -33 411 -27 417
rect -33 399 -27 405
rect -9 411 -3 417
rect -9 399 -3 405
rect 15 411 21 417
rect 15 399 21 405
rect 39 411 45 417
rect 39 399 45 405
rect 63 411 69 417
rect 63 399 69 405
rect 87 411 93 417
rect 87 399 93 405
rect 111 411 117 417
rect 111 399 117 405
rect 135 411 141 417
rect 135 399 141 405
rect 159 411 165 417
rect 159 399 165 405
rect 183 411 189 417
rect 183 399 189 405
rect 207 411 213 417
rect 207 399 213 405
rect 231 411 237 417
rect 231 399 237 405
<< mvpdiffc >>
rect -345 543 -339 549
rect -345 531 -339 537
rect -345 519 -339 525
rect -321 543 -315 549
rect -321 531 -315 537
rect -321 519 -315 525
rect -297 543 -291 549
rect -297 531 -291 537
rect -297 519 -291 525
rect -273 543 -267 549
rect -273 531 -267 537
rect -273 519 -267 525
rect -249 543 -243 549
rect -249 531 -243 537
rect -249 519 -243 525
rect -225 543 -219 549
rect -225 531 -219 537
rect -225 519 -219 525
rect -201 543 -195 549
rect -201 531 -195 537
rect -201 519 -195 525
rect -177 543 -171 549
rect -177 531 -171 537
rect -177 519 -171 525
rect -153 543 -147 549
rect -153 531 -147 537
rect -153 519 -147 525
rect -129 543 -123 549
rect -129 531 -123 537
rect -129 519 -123 525
rect -105 543 -99 549
rect -105 531 -99 537
rect -105 519 -99 525
rect -81 543 -75 549
rect -81 531 -75 537
rect -81 519 -75 525
rect -57 543 -51 549
rect -57 531 -51 537
rect -57 519 -51 525
rect -33 543 -27 549
rect -33 531 -27 537
rect -33 519 -27 525
rect -9 543 -3 549
rect -9 531 -3 537
rect -9 519 -3 525
rect 15 543 21 549
rect 15 531 21 537
rect 15 519 21 525
rect 39 543 45 549
rect 39 531 45 537
rect 39 519 45 525
rect 63 543 69 549
rect 63 531 69 537
rect 63 519 69 525
rect 87 543 93 549
rect 87 531 93 537
rect 87 519 93 525
rect 111 543 117 549
rect 111 531 117 537
rect 111 519 117 525
rect 135 543 141 549
rect 135 531 141 537
rect 135 519 141 525
rect 159 543 165 549
rect 159 531 165 537
rect 159 519 165 525
rect 183 543 189 549
rect 183 531 189 537
rect 183 519 189 525
rect 207 543 213 549
rect 207 531 213 537
rect 207 519 213 525
rect 231 543 237 549
rect 231 531 237 537
rect 231 519 237 525
<< psubdiff >>
rect -396 621 288 624
rect -396 615 -393 621
rect -387 615 -381 621
rect -375 615 -369 621
rect -363 615 -357 621
rect -351 615 -345 621
rect -339 615 -333 621
rect -327 615 -321 621
rect -315 615 -309 621
rect -303 615 -297 621
rect -291 615 -285 621
rect -279 615 -273 621
rect -267 615 -261 621
rect -255 615 -249 621
rect -243 615 -237 621
rect -231 615 -225 621
rect -219 615 -213 621
rect -207 615 -201 621
rect -195 615 -189 621
rect -183 615 -177 621
rect -171 615 -165 621
rect -159 615 -153 621
rect -147 615 -141 621
rect -135 615 -129 621
rect -123 615 -117 621
rect -111 615 -105 621
rect -99 615 -93 621
rect -87 615 -81 621
rect -75 615 -69 621
rect -63 615 -57 621
rect -51 615 -45 621
rect -39 615 -33 621
rect -27 615 -21 621
rect -15 615 -9 621
rect -3 615 3 621
rect 9 615 15 621
rect 21 615 27 621
rect 33 615 39 621
rect 45 615 51 621
rect 57 615 63 621
rect 69 615 75 621
rect 81 615 87 621
rect 93 615 99 621
rect 105 615 111 621
rect 117 615 123 621
rect 129 615 135 621
rect 141 615 147 621
rect 153 615 159 621
rect 165 615 171 621
rect 177 615 183 621
rect 189 615 195 621
rect 201 615 207 621
rect 213 615 219 621
rect 225 615 231 621
rect 237 615 243 621
rect 249 615 255 621
rect 261 615 267 621
rect 273 615 279 621
rect 285 615 288 621
rect -396 612 288 615
rect -396 609 -384 612
rect -396 603 -393 609
rect -387 603 -384 609
rect -396 597 -384 603
rect 276 609 288 612
rect 276 603 279 609
rect 285 603 288 609
rect -396 591 -393 597
rect -387 591 -384 597
rect -396 585 -384 591
rect -396 579 -393 585
rect -387 579 -384 585
rect -396 573 -384 579
rect -396 567 -393 573
rect -387 567 -384 573
rect -396 561 -384 567
rect -396 555 -393 561
rect -387 555 -384 561
rect -396 549 -384 555
rect -396 543 -393 549
rect -387 543 -384 549
rect -396 537 -384 543
rect -396 531 -393 537
rect -387 531 -384 537
rect -396 525 -384 531
rect -396 519 -393 525
rect -387 519 -384 525
rect -396 513 -384 519
rect -396 507 -393 513
rect -387 507 -384 513
rect -396 501 -384 507
rect -396 495 -393 501
rect -387 495 -384 501
rect -396 489 -384 495
rect 276 597 288 603
rect 276 591 279 597
rect 285 591 288 597
rect 276 585 288 591
rect 276 579 279 585
rect 285 579 288 585
rect 276 573 288 579
rect 276 567 279 573
rect 285 567 288 573
rect 276 561 288 567
rect 276 555 279 561
rect 285 555 288 561
rect 276 549 288 555
rect 276 543 279 549
rect 285 543 288 549
rect 276 537 288 543
rect 276 531 279 537
rect 285 531 288 537
rect 276 525 288 531
rect 276 519 279 525
rect 285 519 288 525
rect 276 513 288 519
rect 276 507 279 513
rect 285 507 288 513
rect 276 501 288 507
rect 276 495 279 501
rect 285 495 288 501
rect -396 483 -393 489
rect -387 483 -384 489
rect -396 480 -384 483
rect 276 489 288 495
rect 276 483 279 489
rect 285 483 288 489
rect 276 480 288 483
rect -396 477 288 480
rect -396 471 -393 477
rect -387 471 -381 477
rect -375 471 -369 477
rect -363 471 -357 477
rect -351 471 -345 477
rect -339 471 -333 477
rect -327 471 -321 477
rect -315 471 -309 477
rect -303 471 -297 477
rect -291 471 -285 477
rect -279 471 -273 477
rect -267 471 -261 477
rect -255 471 -249 477
rect -243 471 -237 477
rect -231 471 -225 477
rect -219 471 -213 477
rect -207 471 -201 477
rect -195 471 -189 477
rect -183 471 -177 477
rect -171 471 -165 477
rect -159 471 -153 477
rect -147 471 -141 477
rect -135 471 -129 477
rect -123 471 -117 477
rect -111 471 -105 477
rect -99 471 -93 477
rect -87 471 -81 477
rect -75 471 -69 477
rect -63 471 -57 477
rect -51 471 -45 477
rect -39 471 -33 477
rect -27 471 -21 477
rect -15 471 -9 477
rect -3 471 3 477
rect 9 471 15 477
rect 21 471 27 477
rect 33 471 39 477
rect 45 471 51 477
rect 57 471 63 477
rect 69 471 75 477
rect 81 471 87 477
rect 93 471 99 477
rect 105 471 111 477
rect 117 471 123 477
rect 129 471 135 477
rect 141 471 147 477
rect 153 471 159 477
rect 165 471 171 477
rect 177 471 183 477
rect 189 471 195 477
rect 201 471 207 477
rect 213 471 219 477
rect 225 471 231 477
rect 237 471 243 477
rect 249 471 255 477
rect 261 471 267 477
rect 273 471 279 477
rect 285 471 288 477
rect -396 468 288 471
rect -396 465 -384 468
rect -396 459 -393 465
rect -387 459 -384 465
rect -396 453 -384 459
rect 276 465 288 468
rect 276 459 279 465
rect 285 459 288 465
rect -396 447 -393 453
rect -387 447 -384 453
rect -396 441 -384 447
rect -396 435 -393 441
rect -387 435 -384 441
rect -396 429 -384 435
rect -396 423 -393 429
rect -387 423 -384 429
rect -396 417 -384 423
rect -396 411 -393 417
rect -387 411 -384 417
rect -396 405 -384 411
rect -396 399 -393 405
rect -387 399 -384 405
rect -396 393 -384 399
rect -396 387 -393 393
rect -387 387 -384 393
rect -396 381 -384 387
rect -396 375 -393 381
rect -387 375 -384 381
rect -396 369 -384 375
rect -396 363 -393 369
rect -387 363 -384 369
rect -396 357 -384 363
rect -396 351 -393 357
rect -387 351 -384 357
rect -396 345 -384 351
rect 276 453 288 459
rect 276 447 279 453
rect 285 447 288 453
rect 276 441 288 447
rect 276 435 279 441
rect 285 435 288 441
rect 276 429 288 435
rect 276 423 279 429
rect 285 423 288 429
rect 276 417 288 423
rect 276 411 279 417
rect 285 411 288 417
rect 276 405 288 411
rect 276 399 279 405
rect 285 399 288 405
rect 276 393 288 399
rect 276 387 279 393
rect 285 387 288 393
rect 276 381 288 387
rect 276 375 279 381
rect 285 375 288 381
rect 276 369 288 375
rect 276 363 279 369
rect 285 363 288 369
rect 276 357 288 363
rect 276 351 279 357
rect 285 351 288 357
rect -396 339 -393 345
rect -387 339 -384 345
rect -396 336 -384 339
rect 276 345 288 351
rect 276 339 279 345
rect 285 339 288 345
rect 276 336 288 339
rect -396 333 288 336
rect -396 327 -393 333
rect -387 327 -381 333
rect -375 327 -369 333
rect -363 327 -357 333
rect -351 327 -345 333
rect -339 327 -333 333
rect -327 327 -321 333
rect -315 327 -309 333
rect -303 327 -297 333
rect -291 327 -285 333
rect -279 327 -273 333
rect -267 327 -261 333
rect -255 327 -249 333
rect -243 327 -237 333
rect -231 327 -225 333
rect -219 327 -213 333
rect -207 327 -201 333
rect -195 327 -189 333
rect -183 327 -177 333
rect -171 327 -165 333
rect -159 327 -153 333
rect -147 327 -141 333
rect -135 327 -129 333
rect -123 327 -117 333
rect -111 327 -105 333
rect -99 327 -93 333
rect -87 327 -81 333
rect -75 327 -69 333
rect -63 327 -57 333
rect -51 327 -45 333
rect -39 327 -33 333
rect -27 327 -21 333
rect -15 327 -9 333
rect -3 327 3 333
rect 9 327 15 333
rect 21 327 27 333
rect 33 327 39 333
rect 45 327 51 333
rect 57 327 63 333
rect 69 327 75 333
rect 81 327 87 333
rect 93 327 99 333
rect 105 327 111 333
rect 117 327 123 333
rect 129 327 135 333
rect 141 327 147 333
rect 153 327 159 333
rect 165 327 171 333
rect 177 327 183 333
rect 189 327 195 333
rect 201 327 207 333
rect 213 327 219 333
rect 225 327 231 333
rect 237 327 243 333
rect 249 327 255 333
rect 261 327 267 333
rect 273 327 279 333
rect 285 327 288 333
rect -396 324 288 327
rect -396 321 -384 324
rect -396 315 -393 321
rect -387 315 -384 321
rect -396 309 -384 315
rect -396 303 -393 309
rect -387 303 -384 309
rect -396 297 -384 303
rect -396 291 -393 297
rect -387 291 -384 297
rect -396 285 -384 291
rect -396 279 -393 285
rect -387 279 -384 285
rect -396 273 -384 279
rect -396 267 -393 273
rect -387 267 -384 273
rect -396 261 -384 267
rect -396 255 -393 261
rect -387 255 -384 261
rect -396 249 -384 255
rect -396 243 -393 249
rect -387 243 -384 249
rect -396 237 -384 243
rect -396 231 -393 237
rect -387 231 -384 237
rect -396 225 -384 231
rect -396 219 -393 225
rect -387 219 -384 225
rect -396 213 -384 219
rect -396 207 -393 213
rect -387 207 -384 213
rect -396 201 -384 207
rect -396 195 -393 201
rect -387 195 -384 201
rect -396 189 -384 195
rect -396 183 -393 189
rect -387 183 -384 189
rect -396 177 -384 183
rect -396 171 -393 177
rect -387 171 -384 177
rect -396 165 -384 171
rect -396 159 -393 165
rect -387 159 -384 165
rect -396 153 -384 159
rect -396 147 -393 153
rect -387 147 -384 153
rect -396 141 -384 147
rect -396 135 -393 141
rect -387 135 -384 141
rect -396 129 -384 135
rect -396 123 -393 129
rect -387 123 -384 129
rect -396 117 -384 123
rect -396 111 -393 117
rect -387 111 -384 117
rect -396 105 -384 111
rect -396 99 -393 105
rect -387 99 -384 105
rect -396 96 -384 99
rect 276 321 288 324
rect 276 315 279 321
rect 285 315 288 321
rect 276 309 288 315
rect 276 303 279 309
rect 285 303 288 309
rect 276 297 288 303
rect 276 291 279 297
rect 285 291 288 297
rect 276 285 288 291
rect 276 279 279 285
rect 285 279 288 285
rect 276 273 288 279
rect 276 267 279 273
rect 285 267 288 273
rect 276 261 288 267
rect 276 255 279 261
rect 285 255 288 261
rect 276 249 288 255
rect 276 243 279 249
rect 285 243 288 249
rect 276 237 288 243
rect 276 231 279 237
rect 285 231 288 237
rect 276 225 288 231
rect 276 219 279 225
rect 285 219 288 225
rect 276 213 288 219
rect 276 207 279 213
rect 285 207 288 213
rect 276 201 288 207
rect 276 195 279 201
rect 285 195 288 201
rect 276 189 288 195
rect 276 183 279 189
rect 285 183 288 189
rect 276 177 288 183
rect 276 171 279 177
rect 285 171 288 177
rect 276 165 288 171
rect 276 159 279 165
rect 285 159 288 165
rect 276 153 288 159
rect 276 147 279 153
rect 285 147 288 153
rect 276 141 288 147
rect 276 135 279 141
rect 285 135 288 141
rect 276 129 288 135
rect 276 123 279 129
rect 285 123 288 129
rect 276 117 288 123
rect 276 111 279 117
rect 285 111 288 117
rect 276 105 288 111
rect 276 99 279 105
rect 285 99 288 105
rect 276 96 288 99
rect -396 93 288 96
rect -396 87 -393 93
rect -387 87 -381 93
rect -375 87 -369 93
rect -363 87 -357 93
rect -351 87 -345 93
rect -339 87 -333 93
rect -327 87 -321 93
rect -315 87 -309 93
rect -303 87 -297 93
rect -291 87 -285 93
rect -279 87 -273 93
rect -267 87 -261 93
rect -255 87 -249 93
rect -243 87 -237 93
rect -231 87 -225 93
rect -219 87 -213 93
rect -207 87 -201 93
rect -195 87 -189 93
rect -183 87 -177 93
rect -171 87 -165 93
rect -159 87 -153 93
rect -147 87 -141 93
rect -135 87 -129 93
rect -123 87 -117 93
rect -111 87 -105 93
rect -99 87 -93 93
rect -87 87 -81 93
rect -75 87 -69 93
rect -63 87 -57 93
rect -51 87 -45 93
rect -39 87 -33 93
rect -27 87 -21 93
rect -15 87 -9 93
rect -3 87 3 93
rect 9 87 15 93
rect 21 87 27 93
rect 33 87 39 93
rect 45 87 51 93
rect 57 87 63 93
rect 69 87 75 93
rect 81 87 87 93
rect 93 87 99 93
rect 105 87 111 93
rect 117 87 123 93
rect 129 87 135 93
rect 141 87 147 93
rect 153 87 159 93
rect 165 87 171 93
rect 177 87 183 93
rect 189 87 195 93
rect 201 87 207 93
rect 213 87 219 93
rect 225 87 231 93
rect 237 87 243 93
rect 249 87 255 93
rect 261 87 267 93
rect 273 87 279 93
rect 285 87 288 93
rect -396 84 288 87
rect -396 81 -384 84
rect -396 75 -393 81
rect -387 75 -384 81
rect -396 69 -384 75
rect 276 81 288 84
rect 276 75 279 81
rect 285 75 288 81
rect -396 63 -393 69
rect -387 63 -384 69
rect -396 57 -384 63
rect -396 51 -393 57
rect -387 51 -384 57
rect -396 45 -384 51
rect 276 69 288 75
rect 276 63 279 69
rect 285 63 288 69
rect 276 57 288 63
rect 276 51 279 57
rect 285 51 288 57
rect -396 39 -393 45
rect -387 39 -384 45
rect -396 33 -384 39
rect -396 27 -393 33
rect -387 27 -384 33
rect -396 21 -384 27
rect -396 15 -393 21
rect -387 15 -384 21
rect -396 9 -384 15
rect 276 45 288 51
rect 276 39 279 45
rect 285 39 288 45
rect 276 33 288 39
rect 276 27 279 33
rect 285 27 288 33
rect 276 21 288 27
rect 276 15 279 21
rect 285 15 288 21
rect -396 3 -393 9
rect -387 3 -384 9
rect 276 9 288 15
rect -396 0 -384 3
rect 276 3 279 9
rect 285 3 288 9
rect 276 0 288 3
rect -396 -3 288 0
rect -396 -9 -393 -3
rect -387 -9 -381 -3
rect -375 -9 -369 -3
rect -363 -9 -357 -3
rect -351 -9 -345 -3
rect -339 -9 -333 -3
rect -327 -9 -321 -3
rect -315 -9 -309 -3
rect -303 -9 -297 -3
rect -291 -9 -285 -3
rect -279 -9 -273 -3
rect -267 -9 -261 -3
rect -255 -9 -249 -3
rect -243 -9 -237 -3
rect -231 -9 -225 -3
rect -219 -9 -213 -3
rect -207 -9 -201 -3
rect -195 -9 -189 -3
rect -183 -9 -177 -3
rect -171 -9 -165 -3
rect -159 -9 -153 -3
rect -147 -9 -141 -3
rect -135 -9 -129 -3
rect -123 -9 -117 -3
rect -111 -9 -105 -3
rect -99 -9 -93 -3
rect -87 -9 -81 -3
rect -75 -9 -69 -3
rect -63 -9 -57 -3
rect -51 -9 -45 -3
rect -39 -9 -33 -3
rect -27 -9 -21 -3
rect -15 -9 -9 -3
rect -3 -9 3 -3
rect 9 -9 15 -3
rect 21 -9 27 -3
rect 33 -9 39 -3
rect 45 -9 51 -3
rect 57 -9 63 -3
rect 69 -9 75 -3
rect 81 -9 87 -3
rect 93 -9 99 -3
rect 105 -9 111 -3
rect 117 -9 123 -3
rect 129 -9 135 -3
rect 141 -9 147 -3
rect 153 -9 159 -3
rect 165 -9 171 -3
rect 177 -9 183 -3
rect 189 -9 195 -3
rect 201 -9 207 -3
rect 213 -9 219 -3
rect 225 -9 231 -3
rect 237 -9 243 -3
rect 249 -9 255 -3
rect 261 -9 267 -3
rect 273 -9 279 -3
rect 285 -9 288 -3
rect -396 -12 288 -9
<< nsubdiff >>
rect -372 453 264 456
rect -372 447 -369 453
rect -363 447 -357 453
rect -351 447 -345 453
rect -339 447 -333 453
rect -327 447 -321 453
rect -315 447 -309 453
rect -303 447 -297 453
rect -291 447 -285 453
rect -279 447 -273 453
rect -267 447 -261 453
rect -255 447 -249 453
rect -243 447 -237 453
rect -231 447 -225 453
rect -219 447 -213 453
rect -207 447 -201 453
rect -195 447 -189 453
rect -183 447 -177 453
rect -171 447 -165 453
rect -159 447 -153 453
rect -147 447 -141 453
rect -135 447 -129 453
rect -123 447 -117 453
rect -111 447 -105 453
rect -99 447 -93 453
rect -87 447 -81 453
rect -75 447 -69 453
rect -63 447 -57 453
rect -51 447 -45 453
rect -39 447 -33 453
rect -27 447 -21 453
rect -15 447 -9 453
rect -3 447 3 453
rect 9 447 15 453
rect 21 447 27 453
rect 33 447 39 453
rect 45 447 51 453
rect 57 447 63 453
rect 69 447 75 453
rect 81 447 87 453
rect 93 447 99 453
rect 105 447 111 453
rect 117 447 123 453
rect 129 447 135 453
rect 141 447 147 453
rect 153 447 159 453
rect 165 447 171 453
rect 177 447 183 453
rect 189 447 195 453
rect 201 447 207 453
rect 213 447 219 453
rect 225 447 231 453
rect 237 447 243 453
rect 249 447 255 453
rect 261 447 264 453
rect -372 444 264 447
rect -372 441 -360 444
rect -372 435 -369 441
rect -363 435 -360 441
rect -372 429 -360 435
rect 252 441 264 444
rect 252 435 255 441
rect 261 435 264 441
rect -372 423 -369 429
rect -363 423 -360 429
rect 252 429 264 435
rect -372 417 -360 423
rect -372 411 -369 417
rect -363 411 -360 417
rect -372 405 -360 411
rect -372 399 -369 405
rect -363 399 -360 405
rect -372 393 -360 399
rect 252 423 255 429
rect 261 423 264 429
rect 252 417 264 423
rect 252 411 255 417
rect 261 411 264 417
rect 252 405 264 411
rect 252 399 255 405
rect 261 399 264 405
rect -372 387 -369 393
rect -363 387 -360 393
rect -372 381 -360 387
rect -372 375 -369 381
rect -363 375 -360 381
rect -372 369 -360 375
rect 252 393 264 399
rect 252 387 255 393
rect 261 387 264 393
rect 252 381 264 387
rect 252 375 255 381
rect 261 375 264 381
rect -372 363 -369 369
rect -363 363 -360 369
rect -372 360 -360 363
rect 252 369 264 375
rect 252 363 255 369
rect 261 363 264 369
rect 252 360 264 363
rect -372 357 264 360
rect -372 351 -369 357
rect -363 351 -357 357
rect -351 351 -345 357
rect -339 351 -333 357
rect -327 351 -321 357
rect -315 351 -309 357
rect -303 351 -297 357
rect -291 351 -285 357
rect -279 351 -273 357
rect -267 351 -261 357
rect -255 351 -249 357
rect -243 351 -237 357
rect -231 351 -225 357
rect -219 351 -213 357
rect -207 351 -201 357
rect -195 351 -189 357
rect -183 351 -177 357
rect -171 351 -165 357
rect -159 351 -153 357
rect -147 351 -141 357
rect -135 351 -129 357
rect -123 351 -117 357
rect -111 351 -105 357
rect -99 351 -93 357
rect -87 351 -81 357
rect -75 351 -69 357
rect -63 351 -57 357
rect -51 351 -45 357
rect -39 351 -33 357
rect -27 351 -21 357
rect -15 351 -9 357
rect -3 351 3 357
rect 9 351 15 357
rect 21 351 27 357
rect 33 351 39 357
rect 45 351 51 357
rect 57 351 63 357
rect 69 351 75 357
rect 81 351 87 357
rect 93 351 99 357
rect 105 351 111 357
rect 117 351 123 357
rect 129 351 135 357
rect 141 351 147 357
rect 153 351 159 357
rect 165 351 171 357
rect 177 351 183 357
rect 189 351 195 357
rect 201 351 207 357
rect 213 351 219 357
rect 225 351 231 357
rect 237 351 243 357
rect 249 351 255 357
rect 261 351 264 357
rect -372 348 264 351
<< mvnsubdiff >>
rect -372 597 264 600
rect -372 591 -369 597
rect -363 591 -357 597
rect -351 591 -345 597
rect -339 591 -333 597
rect -327 591 -321 597
rect -315 591 -309 597
rect -303 591 -297 597
rect -291 591 -285 597
rect -279 591 -273 597
rect -267 591 -261 597
rect -255 591 -249 597
rect -243 591 -237 597
rect -231 591 -225 597
rect -219 591 -213 597
rect -207 591 -201 597
rect -195 591 -189 597
rect -183 591 -177 597
rect -171 591 -165 597
rect -159 591 -153 597
rect -147 591 -141 597
rect -135 591 -129 597
rect -123 591 -117 597
rect -111 591 -105 597
rect -99 591 -93 597
rect -87 591 -81 597
rect -75 591 -69 597
rect -63 591 -57 597
rect -51 591 -45 597
rect -39 591 -33 597
rect -27 591 -21 597
rect -15 591 -9 597
rect -3 591 3 597
rect 9 591 15 597
rect 21 591 27 597
rect 33 591 39 597
rect 45 591 51 597
rect 57 591 63 597
rect 69 591 75 597
rect 81 591 87 597
rect 93 591 99 597
rect 105 591 111 597
rect 117 591 123 597
rect 129 591 135 597
rect 141 591 147 597
rect 153 591 159 597
rect 165 591 171 597
rect 177 591 183 597
rect 189 591 195 597
rect 201 591 207 597
rect 213 591 219 597
rect 225 591 231 597
rect 237 591 243 597
rect 249 591 255 597
rect 261 591 264 597
rect -372 588 264 591
rect -372 585 -360 588
rect -372 579 -369 585
rect -363 579 -360 585
rect -372 573 -360 579
rect 252 585 264 588
rect 252 579 255 585
rect 261 579 264 585
rect -372 567 -369 573
rect -363 567 -360 573
rect -372 561 -360 567
rect -372 555 -369 561
rect -363 555 -360 561
rect -372 549 -360 555
rect 252 573 264 579
rect 252 567 255 573
rect 261 567 264 573
rect 252 561 264 567
rect 252 555 255 561
rect 261 555 264 561
rect -372 543 -369 549
rect -363 543 -360 549
rect -372 537 -360 543
rect -372 531 -369 537
rect -363 531 -360 537
rect -372 525 -360 531
rect -372 519 -369 525
rect -363 519 -360 525
rect -372 513 -360 519
rect 252 549 264 555
rect 252 543 255 549
rect 261 543 264 549
rect 252 537 264 543
rect 252 531 255 537
rect 261 531 264 537
rect 252 525 264 531
rect 252 519 255 525
rect 261 519 264 525
rect -372 507 -369 513
rect -363 507 -360 513
rect 252 513 264 519
rect -372 504 -360 507
rect 252 507 255 513
rect 261 507 264 513
rect 252 504 264 507
rect -372 501 264 504
rect -372 495 -369 501
rect -363 495 -357 501
rect -351 495 -345 501
rect -339 495 -333 501
rect -327 495 -321 501
rect -315 495 -309 501
rect -303 495 -297 501
rect -291 495 -285 501
rect -279 495 -273 501
rect -267 495 -261 501
rect -255 495 -249 501
rect -243 495 -237 501
rect -231 495 -225 501
rect -219 495 -213 501
rect -207 495 -201 501
rect -195 495 -189 501
rect -183 495 -177 501
rect -171 495 -165 501
rect -159 495 -153 501
rect -147 495 -141 501
rect -135 495 -129 501
rect -123 495 -117 501
rect -111 495 -105 501
rect -99 495 -93 501
rect -87 495 -81 501
rect -75 495 -69 501
rect -63 495 -57 501
rect -51 495 -45 501
rect -39 495 -33 501
rect -27 495 -21 501
rect -15 495 -9 501
rect -3 495 3 501
rect 9 495 15 501
rect 21 495 27 501
rect 33 495 39 501
rect 45 495 51 501
rect 57 495 63 501
rect 69 495 75 501
rect 81 495 87 501
rect 93 495 99 501
rect 105 495 111 501
rect 117 495 123 501
rect 129 495 135 501
rect 141 495 147 501
rect 153 495 159 501
rect 165 495 171 501
rect 177 495 183 501
rect 189 495 195 501
rect 201 495 207 501
rect 213 495 219 501
rect 225 495 231 501
rect 237 495 243 501
rect 249 495 255 501
rect 261 495 264 501
rect -372 492 264 495
<< psubdiffcont >>
rect -393 615 -387 621
rect -381 615 -375 621
rect -369 615 -363 621
rect -357 615 -351 621
rect -345 615 -339 621
rect -333 615 -327 621
rect -321 615 -315 621
rect -309 615 -303 621
rect -297 615 -291 621
rect -285 615 -279 621
rect -273 615 -267 621
rect -261 615 -255 621
rect -249 615 -243 621
rect -237 615 -231 621
rect -225 615 -219 621
rect -213 615 -207 621
rect -201 615 -195 621
rect -189 615 -183 621
rect -177 615 -171 621
rect -165 615 -159 621
rect -153 615 -147 621
rect -141 615 -135 621
rect -129 615 -123 621
rect -117 615 -111 621
rect -105 615 -99 621
rect -93 615 -87 621
rect -81 615 -75 621
rect -69 615 -63 621
rect -57 615 -51 621
rect -45 615 -39 621
rect -33 615 -27 621
rect -21 615 -15 621
rect -9 615 -3 621
rect 3 615 9 621
rect 15 615 21 621
rect 27 615 33 621
rect 39 615 45 621
rect 51 615 57 621
rect 63 615 69 621
rect 75 615 81 621
rect 87 615 93 621
rect 99 615 105 621
rect 111 615 117 621
rect 123 615 129 621
rect 135 615 141 621
rect 147 615 153 621
rect 159 615 165 621
rect 171 615 177 621
rect 183 615 189 621
rect 195 615 201 621
rect 207 615 213 621
rect 219 615 225 621
rect 231 615 237 621
rect 243 615 249 621
rect 255 615 261 621
rect 267 615 273 621
rect 279 615 285 621
rect -393 603 -387 609
rect 279 603 285 609
rect -393 591 -387 597
rect -393 579 -387 585
rect -393 567 -387 573
rect -393 555 -387 561
rect -393 543 -387 549
rect -393 531 -387 537
rect -393 519 -387 525
rect -393 507 -387 513
rect -393 495 -387 501
rect 279 591 285 597
rect 279 579 285 585
rect 279 567 285 573
rect 279 555 285 561
rect 279 543 285 549
rect 279 531 285 537
rect 279 519 285 525
rect 279 507 285 513
rect 279 495 285 501
rect -393 483 -387 489
rect 279 483 285 489
rect -393 471 -387 477
rect -381 471 -375 477
rect -369 471 -363 477
rect -357 471 -351 477
rect -345 471 -339 477
rect -333 471 -327 477
rect -321 471 -315 477
rect -309 471 -303 477
rect -297 471 -291 477
rect -285 471 -279 477
rect -273 471 -267 477
rect -261 471 -255 477
rect -249 471 -243 477
rect -237 471 -231 477
rect -225 471 -219 477
rect -213 471 -207 477
rect -201 471 -195 477
rect -189 471 -183 477
rect -177 471 -171 477
rect -165 471 -159 477
rect -153 471 -147 477
rect -141 471 -135 477
rect -129 471 -123 477
rect -117 471 -111 477
rect -105 471 -99 477
rect -93 471 -87 477
rect -81 471 -75 477
rect -69 471 -63 477
rect -57 471 -51 477
rect -45 471 -39 477
rect -33 471 -27 477
rect -21 471 -15 477
rect -9 471 -3 477
rect 3 471 9 477
rect 15 471 21 477
rect 27 471 33 477
rect 39 471 45 477
rect 51 471 57 477
rect 63 471 69 477
rect 75 471 81 477
rect 87 471 93 477
rect 99 471 105 477
rect 111 471 117 477
rect 123 471 129 477
rect 135 471 141 477
rect 147 471 153 477
rect 159 471 165 477
rect 171 471 177 477
rect 183 471 189 477
rect 195 471 201 477
rect 207 471 213 477
rect 219 471 225 477
rect 231 471 237 477
rect 243 471 249 477
rect 255 471 261 477
rect 267 471 273 477
rect 279 471 285 477
rect -393 459 -387 465
rect 279 459 285 465
rect -393 447 -387 453
rect -393 435 -387 441
rect -393 423 -387 429
rect -393 411 -387 417
rect -393 399 -387 405
rect -393 387 -387 393
rect -393 375 -387 381
rect -393 363 -387 369
rect -393 351 -387 357
rect 279 447 285 453
rect 279 435 285 441
rect 279 423 285 429
rect 279 411 285 417
rect 279 399 285 405
rect 279 387 285 393
rect 279 375 285 381
rect 279 363 285 369
rect 279 351 285 357
rect -393 339 -387 345
rect 279 339 285 345
rect -393 327 -387 333
rect -381 327 -375 333
rect -369 327 -363 333
rect -357 327 -351 333
rect -345 327 -339 333
rect -333 327 -327 333
rect -321 327 -315 333
rect -309 327 -303 333
rect -297 327 -291 333
rect -285 327 -279 333
rect -273 327 -267 333
rect -261 327 -255 333
rect -249 327 -243 333
rect -237 327 -231 333
rect -225 327 -219 333
rect -213 327 -207 333
rect -201 327 -195 333
rect -189 327 -183 333
rect -177 327 -171 333
rect -165 327 -159 333
rect -153 327 -147 333
rect -141 327 -135 333
rect -129 327 -123 333
rect -117 327 -111 333
rect -105 327 -99 333
rect -93 327 -87 333
rect -81 327 -75 333
rect -69 327 -63 333
rect -57 327 -51 333
rect -45 327 -39 333
rect -33 327 -27 333
rect -21 327 -15 333
rect -9 327 -3 333
rect 3 327 9 333
rect 15 327 21 333
rect 27 327 33 333
rect 39 327 45 333
rect 51 327 57 333
rect 63 327 69 333
rect 75 327 81 333
rect 87 327 93 333
rect 99 327 105 333
rect 111 327 117 333
rect 123 327 129 333
rect 135 327 141 333
rect 147 327 153 333
rect 159 327 165 333
rect 171 327 177 333
rect 183 327 189 333
rect 195 327 201 333
rect 207 327 213 333
rect 219 327 225 333
rect 231 327 237 333
rect 243 327 249 333
rect 255 327 261 333
rect 267 327 273 333
rect 279 327 285 333
rect -393 315 -387 321
rect -393 303 -387 309
rect -393 291 -387 297
rect -393 279 -387 285
rect -393 267 -387 273
rect -393 255 -387 261
rect -393 243 -387 249
rect -393 231 -387 237
rect -393 219 -387 225
rect -393 207 -387 213
rect -393 195 -387 201
rect -393 183 -387 189
rect -393 171 -387 177
rect -393 159 -387 165
rect -393 147 -387 153
rect -393 135 -387 141
rect -393 123 -387 129
rect -393 111 -387 117
rect -393 99 -387 105
rect 279 315 285 321
rect 279 303 285 309
rect 279 291 285 297
rect 279 279 285 285
rect 279 267 285 273
rect 279 255 285 261
rect 279 243 285 249
rect 279 231 285 237
rect 279 219 285 225
rect 279 207 285 213
rect 279 195 285 201
rect 279 183 285 189
rect 279 171 285 177
rect 279 159 285 165
rect 279 147 285 153
rect 279 135 285 141
rect 279 123 285 129
rect 279 111 285 117
rect 279 99 285 105
rect -393 87 -387 93
rect -381 87 -375 93
rect -369 87 -363 93
rect -357 87 -351 93
rect -345 87 -339 93
rect -333 87 -327 93
rect -321 87 -315 93
rect -309 87 -303 93
rect -297 87 -291 93
rect -285 87 -279 93
rect -273 87 -267 93
rect -261 87 -255 93
rect -249 87 -243 93
rect -237 87 -231 93
rect -225 87 -219 93
rect -213 87 -207 93
rect -201 87 -195 93
rect -189 87 -183 93
rect -177 87 -171 93
rect -165 87 -159 93
rect -153 87 -147 93
rect -141 87 -135 93
rect -129 87 -123 93
rect -117 87 -111 93
rect -105 87 -99 93
rect -93 87 -87 93
rect -81 87 -75 93
rect -69 87 -63 93
rect -57 87 -51 93
rect -45 87 -39 93
rect -33 87 -27 93
rect -21 87 -15 93
rect -9 87 -3 93
rect 3 87 9 93
rect 15 87 21 93
rect 27 87 33 93
rect 39 87 45 93
rect 51 87 57 93
rect 63 87 69 93
rect 75 87 81 93
rect 87 87 93 93
rect 99 87 105 93
rect 111 87 117 93
rect 123 87 129 93
rect 135 87 141 93
rect 147 87 153 93
rect 159 87 165 93
rect 171 87 177 93
rect 183 87 189 93
rect 195 87 201 93
rect 207 87 213 93
rect 219 87 225 93
rect 231 87 237 93
rect 243 87 249 93
rect 255 87 261 93
rect 267 87 273 93
rect 279 87 285 93
rect -393 75 -387 81
rect 279 75 285 81
rect -393 63 -387 69
rect -393 51 -387 57
rect 279 63 285 69
rect 279 51 285 57
rect -393 39 -387 45
rect -393 27 -387 33
rect -393 15 -387 21
rect 279 39 285 45
rect 279 27 285 33
rect 279 15 285 21
rect -393 3 -387 9
rect 279 3 285 9
rect -393 -9 -387 -3
rect -381 -9 -375 -3
rect -369 -9 -363 -3
rect -357 -9 -351 -3
rect -345 -9 -339 -3
rect -333 -9 -327 -3
rect -321 -9 -315 -3
rect -309 -9 -303 -3
rect -297 -9 -291 -3
rect -285 -9 -279 -3
rect -273 -9 -267 -3
rect -261 -9 -255 -3
rect -249 -9 -243 -3
rect -237 -9 -231 -3
rect -225 -9 -219 -3
rect -213 -9 -207 -3
rect -201 -9 -195 -3
rect -189 -9 -183 -3
rect -177 -9 -171 -3
rect -165 -9 -159 -3
rect -153 -9 -147 -3
rect -141 -9 -135 -3
rect -129 -9 -123 -3
rect -117 -9 -111 -3
rect -105 -9 -99 -3
rect -93 -9 -87 -3
rect -81 -9 -75 -3
rect -69 -9 -63 -3
rect -57 -9 -51 -3
rect -45 -9 -39 -3
rect -33 -9 -27 -3
rect -21 -9 -15 -3
rect -9 -9 -3 -3
rect 3 -9 9 -3
rect 15 -9 21 -3
rect 27 -9 33 -3
rect 39 -9 45 -3
rect 51 -9 57 -3
rect 63 -9 69 -3
rect 75 -9 81 -3
rect 87 -9 93 -3
rect 99 -9 105 -3
rect 111 -9 117 -3
rect 123 -9 129 -3
rect 135 -9 141 -3
rect 147 -9 153 -3
rect 159 -9 165 -3
rect 171 -9 177 -3
rect 183 -9 189 -3
rect 195 -9 201 -3
rect 207 -9 213 -3
rect 219 -9 225 -3
rect 231 -9 237 -3
rect 243 -9 249 -3
rect 255 -9 261 -3
rect 267 -9 273 -3
rect 279 -9 285 -3
<< nsubdiffcont >>
rect -369 447 -363 453
rect -357 447 -351 453
rect -345 447 -339 453
rect -333 447 -327 453
rect -321 447 -315 453
rect -309 447 -303 453
rect -297 447 -291 453
rect -285 447 -279 453
rect -273 447 -267 453
rect -261 447 -255 453
rect -249 447 -243 453
rect -237 447 -231 453
rect -225 447 -219 453
rect -213 447 -207 453
rect -201 447 -195 453
rect -189 447 -183 453
rect -177 447 -171 453
rect -165 447 -159 453
rect -153 447 -147 453
rect -141 447 -135 453
rect -129 447 -123 453
rect -117 447 -111 453
rect -105 447 -99 453
rect -93 447 -87 453
rect -81 447 -75 453
rect -69 447 -63 453
rect -57 447 -51 453
rect -45 447 -39 453
rect -33 447 -27 453
rect -21 447 -15 453
rect -9 447 -3 453
rect 3 447 9 453
rect 15 447 21 453
rect 27 447 33 453
rect 39 447 45 453
rect 51 447 57 453
rect 63 447 69 453
rect 75 447 81 453
rect 87 447 93 453
rect 99 447 105 453
rect 111 447 117 453
rect 123 447 129 453
rect 135 447 141 453
rect 147 447 153 453
rect 159 447 165 453
rect 171 447 177 453
rect 183 447 189 453
rect 195 447 201 453
rect 207 447 213 453
rect 219 447 225 453
rect 231 447 237 453
rect 243 447 249 453
rect 255 447 261 453
rect -369 435 -363 441
rect 255 435 261 441
rect -369 423 -363 429
rect -369 411 -363 417
rect -369 399 -363 405
rect 255 423 261 429
rect 255 411 261 417
rect 255 399 261 405
rect -369 387 -363 393
rect -369 375 -363 381
rect 255 387 261 393
rect 255 375 261 381
rect -369 363 -363 369
rect 255 363 261 369
rect -369 351 -363 357
rect -357 351 -351 357
rect -345 351 -339 357
rect -333 351 -327 357
rect -321 351 -315 357
rect -309 351 -303 357
rect -297 351 -291 357
rect -285 351 -279 357
rect -273 351 -267 357
rect -261 351 -255 357
rect -249 351 -243 357
rect -237 351 -231 357
rect -225 351 -219 357
rect -213 351 -207 357
rect -201 351 -195 357
rect -189 351 -183 357
rect -177 351 -171 357
rect -165 351 -159 357
rect -153 351 -147 357
rect -141 351 -135 357
rect -129 351 -123 357
rect -117 351 -111 357
rect -105 351 -99 357
rect -93 351 -87 357
rect -81 351 -75 357
rect -69 351 -63 357
rect -57 351 -51 357
rect -45 351 -39 357
rect -33 351 -27 357
rect -21 351 -15 357
rect -9 351 -3 357
rect 3 351 9 357
rect 15 351 21 357
rect 27 351 33 357
rect 39 351 45 357
rect 51 351 57 357
rect 63 351 69 357
rect 75 351 81 357
rect 87 351 93 357
rect 99 351 105 357
rect 111 351 117 357
rect 123 351 129 357
rect 135 351 141 357
rect 147 351 153 357
rect 159 351 165 357
rect 171 351 177 357
rect 183 351 189 357
rect 195 351 201 357
rect 207 351 213 357
rect 219 351 225 357
rect 231 351 237 357
rect 243 351 249 357
rect 255 351 261 357
<< mvnsubdiffcont >>
rect -369 591 -363 597
rect -357 591 -351 597
rect -345 591 -339 597
rect -333 591 -327 597
rect -321 591 -315 597
rect -309 591 -303 597
rect -297 591 -291 597
rect -285 591 -279 597
rect -273 591 -267 597
rect -261 591 -255 597
rect -249 591 -243 597
rect -237 591 -231 597
rect -225 591 -219 597
rect -213 591 -207 597
rect -201 591 -195 597
rect -189 591 -183 597
rect -177 591 -171 597
rect -165 591 -159 597
rect -153 591 -147 597
rect -141 591 -135 597
rect -129 591 -123 597
rect -117 591 -111 597
rect -105 591 -99 597
rect -93 591 -87 597
rect -81 591 -75 597
rect -69 591 -63 597
rect -57 591 -51 597
rect -45 591 -39 597
rect -33 591 -27 597
rect -21 591 -15 597
rect -9 591 -3 597
rect 3 591 9 597
rect 15 591 21 597
rect 27 591 33 597
rect 39 591 45 597
rect 51 591 57 597
rect 63 591 69 597
rect 75 591 81 597
rect 87 591 93 597
rect 99 591 105 597
rect 111 591 117 597
rect 123 591 129 597
rect 135 591 141 597
rect 147 591 153 597
rect 159 591 165 597
rect 171 591 177 597
rect 183 591 189 597
rect 195 591 201 597
rect 207 591 213 597
rect 219 591 225 597
rect 231 591 237 597
rect 243 591 249 597
rect 255 591 261 597
rect -369 579 -363 585
rect 255 579 261 585
rect -369 567 -363 573
rect -369 555 -363 561
rect 255 567 261 573
rect 255 555 261 561
rect -369 543 -363 549
rect -369 531 -363 537
rect -369 519 -363 525
rect 255 543 261 549
rect 255 531 261 537
rect 255 519 261 525
rect -369 507 -363 513
rect 255 507 261 513
rect -369 495 -363 501
rect -357 495 -351 501
rect -345 495 -339 501
rect -333 495 -327 501
rect -321 495 -315 501
rect -309 495 -303 501
rect -297 495 -291 501
rect -285 495 -279 501
rect -273 495 -267 501
rect -261 495 -255 501
rect -249 495 -243 501
rect -237 495 -231 501
rect -225 495 -219 501
rect -213 495 -207 501
rect -201 495 -195 501
rect -189 495 -183 501
rect -177 495 -171 501
rect -165 495 -159 501
rect -153 495 -147 501
rect -141 495 -135 501
rect -129 495 -123 501
rect -117 495 -111 501
rect -105 495 -99 501
rect -93 495 -87 501
rect -81 495 -75 501
rect -69 495 -63 501
rect -57 495 -51 501
rect -45 495 -39 501
rect -33 495 -27 501
rect -21 495 -15 501
rect -9 495 -3 501
rect 3 495 9 501
rect 15 495 21 501
rect 27 495 33 501
rect 39 495 45 501
rect 51 495 57 501
rect 63 495 69 501
rect 75 495 81 501
rect 87 495 93 501
rect 99 495 105 501
rect 111 495 117 501
rect 123 495 129 501
rect 135 495 141 501
rect 147 495 153 501
rect 159 495 165 501
rect 171 495 177 501
rect 183 495 189 501
rect 195 495 201 501
rect 207 495 213 501
rect 219 495 225 501
rect 231 495 237 501
rect 243 495 249 501
rect 255 495 261 501
<< polysilicon >>
rect -336 573 -300 576
rect -336 567 -333 573
rect -327 567 -321 573
rect -315 567 -309 573
rect -303 567 -300 573
rect -336 564 -300 567
rect -336 552 -324 564
rect -312 552 -300 564
rect -288 573 -252 576
rect -288 567 -285 573
rect -279 567 -273 573
rect -267 567 -261 573
rect -255 567 -252 573
rect -288 564 -252 567
rect -288 552 -276 564
rect -264 552 -252 564
rect -240 573 -204 576
rect -240 567 -237 573
rect -231 567 -225 573
rect -219 567 -213 573
rect -207 567 -204 573
rect -240 564 -204 567
rect -240 552 -228 564
rect -216 552 -204 564
rect -192 573 -156 576
rect -192 567 -189 573
rect -183 567 -177 573
rect -171 567 -165 573
rect -159 567 -156 573
rect -192 564 -156 567
rect -192 552 -180 564
rect -168 552 -156 564
rect -144 573 -108 576
rect -144 567 -141 573
rect -135 567 -129 573
rect -123 567 -117 573
rect -111 567 -108 573
rect -144 564 -108 567
rect -144 552 -132 564
rect -120 552 -108 564
rect -96 573 -60 576
rect -96 567 -93 573
rect -87 567 -81 573
rect -75 567 -69 573
rect -63 567 -60 573
rect -96 564 -60 567
rect -96 552 -84 564
rect -72 552 -60 564
rect -48 573 -12 576
rect -48 567 -45 573
rect -39 567 -33 573
rect -27 567 -21 573
rect -15 567 -12 573
rect -48 564 -12 567
rect -48 552 -36 564
rect -24 552 -12 564
rect 0 573 36 576
rect 0 567 3 573
rect 9 567 15 573
rect 21 567 27 573
rect 33 567 36 573
rect 0 564 36 567
rect 0 552 12 564
rect 24 552 36 564
rect 48 573 84 576
rect 48 567 51 573
rect 57 567 63 573
rect 69 567 75 573
rect 81 567 84 573
rect 48 564 84 567
rect 48 552 60 564
rect 72 552 84 564
rect 96 573 132 576
rect 96 567 99 573
rect 105 567 111 573
rect 117 567 123 573
rect 129 567 132 573
rect 96 564 132 567
rect 96 552 108 564
rect 120 552 132 564
rect 144 573 180 576
rect 144 567 147 573
rect 153 567 159 573
rect 165 567 171 573
rect 177 567 180 573
rect 144 564 180 567
rect 144 552 156 564
rect 168 552 180 564
rect 192 573 228 576
rect 192 567 195 573
rect 201 567 207 573
rect 213 567 219 573
rect 225 567 228 573
rect 192 564 228 567
rect 192 552 204 564
rect 216 552 228 564
rect -336 510 -324 516
rect -312 510 -300 516
rect -288 510 -276 516
rect -264 510 -252 516
rect -240 510 -228 516
rect -216 510 -204 516
rect -192 510 -180 516
rect -168 510 -156 516
rect -144 510 -132 516
rect -120 510 -108 516
rect -96 510 -84 516
rect -72 510 -60 516
rect -48 510 -36 516
rect -24 510 -12 516
rect 0 510 12 516
rect 24 510 36 516
rect 48 510 60 516
rect 72 510 84 516
rect 96 510 108 516
rect 120 510 132 516
rect 144 510 156 516
rect 168 510 180 516
rect 192 510 204 516
rect 216 510 228 516
rect -336 426 -324 432
rect -312 426 -300 432
rect -288 426 -276 432
rect -264 426 -252 432
rect -240 426 -228 432
rect -216 426 -204 432
rect -192 426 -180 432
rect -168 426 -156 432
rect -144 426 -132 432
rect -120 426 -108 432
rect -96 426 -84 432
rect -72 426 -60 432
rect -48 426 -36 432
rect -24 426 -12 432
rect 0 426 12 432
rect 24 426 36 432
rect 48 426 60 432
rect 72 426 84 432
rect 96 426 108 432
rect 120 426 132 432
rect 144 426 156 432
rect 168 426 180 432
rect 192 426 204 432
rect 216 426 228 432
rect -336 384 -324 396
rect -312 384 -300 396
rect -336 381 -300 384
rect -336 375 -333 381
rect -327 375 -321 381
rect -315 375 -309 381
rect -303 375 -300 381
rect -336 372 -300 375
rect -288 384 -276 396
rect -264 384 -252 396
rect -288 381 -252 384
rect -288 375 -285 381
rect -279 375 -273 381
rect -267 375 -261 381
rect -255 375 -252 381
rect -288 372 -252 375
rect -240 384 -228 396
rect -216 384 -204 396
rect -240 381 -204 384
rect -240 375 -237 381
rect -231 375 -225 381
rect -219 375 -213 381
rect -207 375 -204 381
rect -240 372 -204 375
rect -192 384 -180 396
rect -168 384 -156 396
rect -192 381 -156 384
rect -192 375 -189 381
rect -183 375 -177 381
rect -171 375 -165 381
rect -159 375 -156 381
rect -192 372 -156 375
rect -144 384 -132 396
rect -120 384 -108 396
rect -144 381 -108 384
rect -144 375 -141 381
rect -135 375 -129 381
rect -123 375 -117 381
rect -111 375 -108 381
rect -144 372 -108 375
rect -96 384 -84 396
rect -72 384 -60 396
rect -96 381 -60 384
rect -96 375 -93 381
rect -87 375 -81 381
rect -75 375 -69 381
rect -63 375 -60 381
rect -96 372 -60 375
rect -48 384 -36 396
rect -24 384 -12 396
rect -48 381 -12 384
rect -48 375 -45 381
rect -39 375 -33 381
rect -27 375 -21 381
rect -15 375 -12 381
rect -48 372 -12 375
rect 0 384 12 396
rect 24 384 36 396
rect 0 381 36 384
rect 0 375 3 381
rect 9 375 15 381
rect 21 375 27 381
rect 33 375 36 381
rect 0 372 36 375
rect 48 384 60 396
rect 72 384 84 396
rect 48 381 84 384
rect 48 375 51 381
rect 57 375 63 381
rect 69 375 75 381
rect 81 375 84 381
rect 48 372 84 375
rect 96 384 108 396
rect 120 384 132 396
rect 96 381 132 384
rect 96 375 99 381
rect 105 375 111 381
rect 117 375 123 381
rect 129 375 132 381
rect 96 372 132 375
rect 144 384 156 396
rect 168 384 180 396
rect 144 381 180 384
rect 144 375 147 381
rect 153 375 159 381
rect 165 375 171 381
rect 177 375 180 381
rect 144 372 180 375
rect 192 384 204 396
rect 216 384 228 396
rect 192 381 228 384
rect 192 375 195 381
rect 201 375 207 381
rect 213 375 219 381
rect 225 375 228 381
rect 192 372 228 375
rect -336 69 -300 72
rect -336 63 -333 69
rect -327 63 -321 69
rect -315 63 -309 69
rect -303 63 -300 69
rect -336 60 -300 63
rect -336 48 -324 60
rect -312 48 -300 60
rect -288 69 -252 72
rect -288 63 -285 69
rect -279 63 -273 69
rect -267 63 -261 69
rect -255 63 -252 69
rect -288 60 -252 63
rect -288 48 -276 60
rect -264 48 -252 60
rect -240 69 -204 72
rect -240 63 -237 69
rect -231 63 -225 69
rect -219 63 -213 69
rect -207 63 -204 69
rect -240 60 -204 63
rect -240 48 -228 60
rect -216 48 -204 60
rect -192 69 -156 72
rect -192 63 -189 69
rect -183 63 -177 69
rect -171 63 -165 69
rect -159 63 -156 69
rect -192 60 -156 63
rect -192 48 -180 60
rect -168 48 -156 60
rect -144 69 -108 72
rect -144 63 -141 69
rect -135 63 -129 69
rect -123 63 -117 69
rect -111 63 -108 69
rect -144 60 -108 63
rect -144 48 -132 60
rect -120 48 -108 60
rect -96 69 -60 72
rect -96 63 -93 69
rect -87 63 -81 69
rect -75 63 -69 69
rect -63 63 -60 69
rect -96 60 -60 63
rect -96 48 -84 60
rect -72 48 -60 60
rect -48 69 -12 72
rect -48 63 -45 69
rect -39 63 -33 69
rect -27 63 -21 69
rect -15 63 -12 69
rect -48 60 -12 63
rect -48 48 -36 60
rect -24 48 -12 60
rect 0 69 36 72
rect 0 63 3 69
rect 9 63 15 69
rect 21 63 27 69
rect 33 63 36 69
rect 0 60 36 63
rect 0 48 12 60
rect 24 48 36 60
rect 48 69 84 72
rect 48 63 51 69
rect 57 63 63 69
rect 69 63 75 69
rect 81 63 84 69
rect 48 60 84 63
rect 48 48 60 60
rect 72 48 84 60
rect 96 69 132 72
rect 96 63 99 69
rect 105 63 111 69
rect 117 63 123 69
rect 129 63 132 69
rect 96 60 132 63
rect 96 48 108 60
rect 120 48 132 60
rect 144 69 180 72
rect 144 63 147 69
rect 153 63 159 69
rect 165 63 171 69
rect 177 63 180 69
rect 144 60 180 63
rect 144 48 156 60
rect 168 48 180 60
rect 192 69 228 72
rect 192 63 195 69
rect 201 63 207 69
rect 213 63 219 69
rect 225 63 228 69
rect 192 60 228 63
rect 192 48 204 60
rect 216 48 228 60
rect -336 6 -324 12
rect -312 6 -300 12
rect -288 6 -276 12
rect -264 6 -252 12
rect -240 6 -228 12
rect -216 6 -204 12
rect -192 6 -180 12
rect -168 6 -156 12
rect -144 6 -132 12
rect -120 6 -108 12
rect -96 6 -84 12
rect -72 6 -60 12
rect -48 6 -36 12
rect -24 6 -12 12
rect 0 6 12 12
rect 24 6 36 12
rect 48 6 60 12
rect 72 6 84 12
rect 96 6 108 12
rect 120 6 132 12
rect 144 6 156 12
rect 168 6 180 12
rect 192 6 204 12
rect 216 6 228 12
<< polycontact >>
rect -333 567 -327 573
rect -321 567 -315 573
rect -309 567 -303 573
rect -285 567 -279 573
rect -273 567 -267 573
rect -261 567 -255 573
rect -237 567 -231 573
rect -225 567 -219 573
rect -213 567 -207 573
rect -189 567 -183 573
rect -177 567 -171 573
rect -165 567 -159 573
rect -141 567 -135 573
rect -129 567 -123 573
rect -117 567 -111 573
rect -93 567 -87 573
rect -81 567 -75 573
rect -69 567 -63 573
rect -45 567 -39 573
rect -33 567 -27 573
rect -21 567 -15 573
rect 3 567 9 573
rect 15 567 21 573
rect 27 567 33 573
rect 51 567 57 573
rect 63 567 69 573
rect 75 567 81 573
rect 99 567 105 573
rect 111 567 117 573
rect 123 567 129 573
rect 147 567 153 573
rect 159 567 165 573
rect 171 567 177 573
rect 195 567 201 573
rect 207 567 213 573
rect 219 567 225 573
rect -333 375 -327 381
rect -321 375 -315 381
rect -309 375 -303 381
rect -285 375 -279 381
rect -273 375 -267 381
rect -261 375 -255 381
rect -237 375 -231 381
rect -225 375 -219 381
rect -213 375 -207 381
rect -189 375 -183 381
rect -177 375 -171 381
rect -165 375 -159 381
rect -141 375 -135 381
rect -129 375 -123 381
rect -117 375 -111 381
rect -93 375 -87 381
rect -81 375 -75 381
rect -69 375 -63 381
rect -45 375 -39 381
rect -33 375 -27 381
rect -21 375 -15 381
rect 3 375 9 381
rect 15 375 21 381
rect 27 375 33 381
rect 51 375 57 381
rect 63 375 69 381
rect 75 375 81 381
rect 99 375 105 381
rect 111 375 117 381
rect 123 375 129 381
rect 147 375 153 381
rect 159 375 165 381
rect 171 375 177 381
rect 195 375 201 381
rect 207 375 213 381
rect 219 375 225 381
rect -333 63 -327 69
rect -321 63 -315 69
rect -309 63 -303 69
rect -285 63 -279 69
rect -273 63 -267 69
rect -261 63 -255 69
rect -237 63 -231 69
rect -225 63 -219 69
rect -213 63 -207 69
rect -189 63 -183 69
rect -177 63 -171 69
rect -165 63 -159 69
rect -141 63 -135 69
rect -129 63 -123 69
rect -117 63 -111 69
rect -93 63 -87 69
rect -81 63 -75 69
rect -69 63 -63 69
rect -45 63 -39 69
rect -33 63 -27 69
rect -21 63 -15 69
rect 3 63 9 69
rect 15 63 21 69
rect 27 63 33 69
rect 51 63 57 69
rect 63 63 69 69
rect 75 63 81 69
rect 99 63 105 69
rect 111 63 117 69
rect 123 63 129 69
rect 147 63 153 69
rect 159 63 165 69
rect 171 63 177 69
rect 195 63 201 69
rect 207 63 213 69
rect 219 63 225 69
<< metal1 >>
rect -396 621 288 624
rect -396 615 -393 621
rect -387 615 -381 621
rect -375 615 -369 621
rect -363 615 -357 621
rect -351 615 -345 621
rect -339 615 -333 621
rect -327 615 -321 621
rect -315 615 -309 621
rect -303 615 -297 621
rect -291 615 -285 621
rect -279 615 -273 621
rect -267 615 -261 621
rect -255 615 -249 621
rect -243 615 -237 621
rect -231 615 -225 621
rect -219 615 -213 621
rect -207 615 -201 621
rect -195 615 -189 621
rect -183 615 -177 621
rect -171 615 -165 621
rect -159 615 -153 621
rect -147 615 -141 621
rect -135 615 -129 621
rect -123 615 -117 621
rect -111 615 -105 621
rect -99 615 -93 621
rect -87 615 -81 621
rect -75 615 -69 621
rect -63 615 -57 621
rect -51 615 -45 621
rect -39 615 -33 621
rect -27 615 -21 621
rect -15 615 -9 621
rect -3 615 3 621
rect 9 615 15 621
rect 21 615 27 621
rect 33 615 39 621
rect 45 615 51 621
rect 57 615 63 621
rect 69 615 75 621
rect 81 615 87 621
rect 93 615 99 621
rect 105 615 111 621
rect 117 615 123 621
rect 129 615 135 621
rect 141 615 147 621
rect 153 615 159 621
rect 165 615 171 621
rect 177 615 183 621
rect 189 615 195 621
rect 201 615 207 621
rect 213 615 219 621
rect 225 615 231 621
rect 237 615 243 621
rect 249 615 255 621
rect 261 615 267 621
rect 273 615 279 621
rect 285 615 288 621
rect -396 612 288 615
rect -396 609 -384 612
rect -396 603 -393 609
rect -387 603 -384 609
rect -396 597 -384 603
rect 276 609 288 612
rect 276 603 279 609
rect 285 603 288 609
rect -396 591 -393 597
rect -387 591 -384 597
rect -396 585 -384 591
rect -396 579 -393 585
rect -387 579 -384 585
rect -396 573 -384 579
rect -396 567 -393 573
rect -387 567 -384 573
rect -396 561 -384 567
rect -396 555 -393 561
rect -387 555 -384 561
rect -396 549 -384 555
rect -396 543 -393 549
rect -387 543 -384 549
rect -396 537 -384 543
rect -396 531 -393 537
rect -387 531 -384 537
rect -396 525 -384 531
rect -396 519 -393 525
rect -387 519 -384 525
rect -396 513 -384 519
rect -396 507 -393 513
rect -387 507 -384 513
rect -396 501 -384 507
rect -396 495 -393 501
rect -387 495 -384 501
rect -396 489 -384 495
rect -372 597 264 600
rect -372 591 -369 597
rect -363 591 -357 597
rect -351 591 -345 597
rect -339 591 -333 597
rect -327 591 -321 597
rect -315 591 -309 597
rect -303 591 -297 597
rect -291 591 -285 597
rect -279 591 -273 597
rect -267 591 -261 597
rect -255 591 -249 597
rect -243 591 -237 597
rect -231 591 -225 597
rect -219 591 -213 597
rect -207 591 -201 597
rect -195 591 -189 597
rect -183 591 -177 597
rect -171 591 -165 597
rect -159 591 -153 597
rect -147 591 -141 597
rect -135 591 -129 597
rect -123 591 -117 597
rect -111 591 -105 597
rect -99 591 -93 597
rect -87 591 -81 597
rect -75 591 -69 597
rect -63 591 -57 597
rect -51 591 -45 597
rect -39 591 -33 597
rect -27 591 -21 597
rect -15 591 -9 597
rect -3 591 3 597
rect 9 591 15 597
rect 21 591 27 597
rect 33 591 39 597
rect 45 591 51 597
rect 57 591 63 597
rect 69 591 75 597
rect 81 591 87 597
rect 93 591 99 597
rect 105 591 111 597
rect 117 591 123 597
rect 129 591 135 597
rect 141 591 147 597
rect 153 591 159 597
rect 165 591 171 597
rect 177 591 183 597
rect 189 591 195 597
rect 201 591 207 597
rect 213 591 219 597
rect 225 591 231 597
rect 237 591 243 597
rect 249 591 255 597
rect 261 591 264 597
rect -372 588 264 591
rect -372 585 -360 588
rect -372 579 -369 585
rect -363 579 -360 585
rect -372 573 -360 579
rect 252 585 264 588
rect 252 579 255 585
rect 261 579 264 585
rect -372 567 -369 573
rect -363 567 -360 573
rect -372 561 -360 567
rect -336 573 -300 576
rect -336 567 -333 573
rect -327 567 -321 573
rect -315 567 -309 573
rect -303 567 -300 573
rect -336 564 -300 567
rect -288 573 -252 576
rect -288 567 -285 573
rect -279 567 -273 573
rect -267 567 -261 573
rect -255 567 -252 573
rect -288 564 -252 567
rect -240 573 -204 576
rect -240 567 -237 573
rect -231 567 -225 573
rect -219 567 -213 573
rect -207 567 -204 573
rect -240 564 -204 567
rect -192 573 -156 576
rect -192 567 -189 573
rect -183 567 -177 573
rect -171 567 -165 573
rect -159 567 -156 573
rect -192 564 -156 567
rect -144 573 -108 576
rect -144 567 -141 573
rect -135 567 -129 573
rect -123 567 -117 573
rect -111 567 -108 573
rect -144 564 -108 567
rect -96 573 -60 576
rect -96 567 -93 573
rect -87 567 -81 573
rect -75 567 -69 573
rect -63 567 -60 573
rect -96 564 -60 567
rect -48 573 -12 576
rect -48 567 -45 573
rect -39 567 -33 573
rect -27 567 -21 573
rect -15 567 -12 573
rect -48 564 -12 567
rect 0 573 36 576
rect 0 567 3 573
rect 9 567 15 573
rect 21 567 27 573
rect 33 567 36 573
rect 0 564 36 567
rect 48 573 84 576
rect 48 567 51 573
rect 57 567 63 573
rect 69 567 75 573
rect 81 567 84 573
rect 48 564 84 567
rect 96 573 132 576
rect 96 567 99 573
rect 105 567 111 573
rect 117 567 123 573
rect 129 567 132 573
rect 96 564 132 567
rect 144 573 180 576
rect 144 567 147 573
rect 153 567 159 573
rect 165 567 171 573
rect 177 567 180 573
rect 144 564 180 567
rect 192 573 228 576
rect 192 567 195 573
rect 201 567 207 573
rect 213 567 219 573
rect 225 567 228 573
rect 192 564 228 567
rect 252 573 264 579
rect 252 567 255 573
rect 261 567 264 573
rect -372 555 -369 561
rect -363 555 -360 561
rect -372 549 -360 555
rect 252 561 264 567
rect 252 555 255 561
rect 261 555 264 561
rect -372 543 -369 549
rect -363 543 -360 549
rect -372 537 -360 543
rect -372 531 -369 537
rect -363 531 -360 537
rect -372 525 -360 531
rect -372 519 -369 525
rect -363 519 -360 525
rect -372 513 -360 519
rect -372 507 -369 513
rect -363 507 -360 513
rect -372 504 -360 507
rect -348 549 -336 552
rect -348 543 -345 549
rect -339 543 -336 549
rect -348 537 -336 543
rect -348 531 -345 537
rect -339 531 -336 537
rect -348 525 -336 531
rect -348 519 -345 525
rect -339 519 -336 525
rect -348 504 -336 519
rect -324 549 -312 552
rect -324 543 -321 549
rect -315 543 -312 549
rect -324 537 -312 543
rect -324 531 -321 537
rect -315 531 -312 537
rect -324 525 -312 531
rect -324 519 -321 525
rect -315 519 -312 525
rect -324 516 -312 519
rect -300 549 -288 552
rect -300 543 -297 549
rect -291 543 -288 549
rect -300 537 -288 543
rect -300 531 -297 537
rect -291 531 -288 537
rect -300 525 -288 531
rect -300 519 -297 525
rect -291 519 -288 525
rect -300 504 -288 519
rect -276 549 -264 552
rect -276 543 -273 549
rect -267 543 -264 549
rect -276 537 -264 543
rect -276 531 -273 537
rect -267 531 -264 537
rect -276 525 -264 531
rect -276 519 -273 525
rect -267 519 -264 525
rect -276 516 -264 519
rect -252 549 -240 552
rect -252 543 -249 549
rect -243 543 -240 549
rect -252 537 -240 543
rect -252 531 -249 537
rect -243 531 -240 537
rect -252 525 -240 531
rect -252 519 -249 525
rect -243 519 -240 525
rect -252 504 -240 519
rect -228 549 -216 552
rect -228 543 -225 549
rect -219 543 -216 549
rect -228 537 -216 543
rect -228 531 -225 537
rect -219 531 -216 537
rect -228 525 -216 531
rect -228 519 -225 525
rect -219 519 -216 525
rect -228 516 -216 519
rect -204 549 -192 552
rect -204 543 -201 549
rect -195 543 -192 549
rect -204 537 -192 543
rect -204 531 -201 537
rect -195 531 -192 537
rect -204 525 -192 531
rect -204 519 -201 525
rect -195 519 -192 525
rect -204 504 -192 519
rect -180 549 -168 552
rect -180 543 -177 549
rect -171 543 -168 549
rect -180 537 -168 543
rect -180 531 -177 537
rect -171 531 -168 537
rect -180 525 -168 531
rect -180 519 -177 525
rect -171 519 -168 525
rect -180 516 -168 519
rect -156 549 -144 552
rect -156 543 -153 549
rect -147 543 -144 549
rect -156 537 -144 543
rect -156 531 -153 537
rect -147 531 -144 537
rect -156 525 -144 531
rect -156 519 -153 525
rect -147 519 -144 525
rect -156 504 -144 519
rect -132 549 -120 552
rect -132 543 -129 549
rect -123 543 -120 549
rect -132 537 -120 543
rect -132 531 -129 537
rect -123 531 -120 537
rect -132 525 -120 531
rect -132 519 -129 525
rect -123 519 -120 525
rect -132 516 -120 519
rect -108 549 -96 552
rect -108 543 -105 549
rect -99 543 -96 549
rect -108 537 -96 543
rect -108 531 -105 537
rect -99 531 -96 537
rect -108 525 -96 531
rect -108 519 -105 525
rect -99 519 -96 525
rect -108 504 -96 519
rect -84 549 -72 552
rect -84 543 -81 549
rect -75 543 -72 549
rect -84 537 -72 543
rect -84 531 -81 537
rect -75 531 -72 537
rect -84 525 -72 531
rect -84 519 -81 525
rect -75 519 -72 525
rect -84 516 -72 519
rect -60 549 -48 552
rect -60 543 -57 549
rect -51 543 -48 549
rect -60 537 -48 543
rect -60 531 -57 537
rect -51 531 -48 537
rect -60 525 -48 531
rect -60 519 -57 525
rect -51 519 -48 525
rect -60 504 -48 519
rect -36 549 -24 552
rect -36 543 -33 549
rect -27 543 -24 549
rect -36 537 -24 543
rect -36 531 -33 537
rect -27 531 -24 537
rect -36 525 -24 531
rect -36 519 -33 525
rect -27 519 -24 525
rect -36 516 -24 519
rect -12 549 0 552
rect -12 543 -9 549
rect -3 543 0 549
rect -12 537 0 543
rect -12 531 -9 537
rect -3 531 0 537
rect -12 525 0 531
rect -12 519 -9 525
rect -3 519 0 525
rect -12 504 0 519
rect 12 549 24 552
rect 12 543 15 549
rect 21 543 24 549
rect 12 537 24 543
rect 12 531 15 537
rect 21 531 24 537
rect 12 525 24 531
rect 12 519 15 525
rect 21 519 24 525
rect 12 516 24 519
rect 36 549 48 552
rect 36 543 39 549
rect 45 543 48 549
rect 36 537 48 543
rect 36 531 39 537
rect 45 531 48 537
rect 36 525 48 531
rect 36 519 39 525
rect 45 519 48 525
rect 36 504 48 519
rect 60 549 72 552
rect 60 543 63 549
rect 69 543 72 549
rect 60 537 72 543
rect 60 531 63 537
rect 69 531 72 537
rect 60 525 72 531
rect 60 519 63 525
rect 69 519 72 525
rect 60 516 72 519
rect 84 549 96 552
rect 84 543 87 549
rect 93 543 96 549
rect 84 537 96 543
rect 84 531 87 537
rect 93 531 96 537
rect 84 525 96 531
rect 84 519 87 525
rect 93 519 96 525
rect 84 504 96 519
rect 108 549 120 552
rect 108 543 111 549
rect 117 543 120 549
rect 108 537 120 543
rect 108 531 111 537
rect 117 531 120 537
rect 108 525 120 531
rect 108 519 111 525
rect 117 519 120 525
rect 108 516 120 519
rect 132 549 144 552
rect 132 543 135 549
rect 141 543 144 549
rect 132 537 144 543
rect 132 531 135 537
rect 141 531 144 537
rect 132 525 144 531
rect 132 519 135 525
rect 141 519 144 525
rect 132 504 144 519
rect 156 549 168 552
rect 156 543 159 549
rect 165 543 168 549
rect 156 537 168 543
rect 156 531 159 537
rect 165 531 168 537
rect 156 525 168 531
rect 156 519 159 525
rect 165 519 168 525
rect 156 516 168 519
rect 180 549 192 552
rect 180 543 183 549
rect 189 543 192 549
rect 180 537 192 543
rect 180 531 183 537
rect 189 531 192 537
rect 180 525 192 531
rect 180 519 183 525
rect 189 519 192 525
rect 180 504 192 519
rect 204 549 216 552
rect 204 543 207 549
rect 213 543 216 549
rect 204 537 216 543
rect 204 531 207 537
rect 213 531 216 537
rect 204 525 216 531
rect 204 519 207 525
rect 213 519 216 525
rect 204 516 216 519
rect 228 549 240 552
rect 228 543 231 549
rect 237 543 240 549
rect 228 537 240 543
rect 228 531 231 537
rect 237 531 240 537
rect 228 525 240 531
rect 228 519 231 525
rect 237 519 240 525
rect 228 504 240 519
rect 252 549 264 555
rect 252 543 255 549
rect 261 543 264 549
rect 252 537 264 543
rect 252 531 255 537
rect 261 531 264 537
rect 252 525 264 531
rect 252 519 255 525
rect 261 519 264 525
rect 252 513 264 519
rect 252 507 255 513
rect 261 507 264 513
rect 252 504 264 507
rect -372 501 264 504
rect -372 495 -369 501
rect -363 495 -357 501
rect -351 495 -345 501
rect -339 495 -333 501
rect -327 495 -321 501
rect -315 495 -309 501
rect -303 495 -297 501
rect -291 495 -285 501
rect -279 495 -273 501
rect -267 495 -261 501
rect -255 495 -249 501
rect -243 495 -237 501
rect -231 495 -225 501
rect -219 495 -213 501
rect -207 495 -201 501
rect -195 495 -189 501
rect -183 495 -177 501
rect -171 495 -165 501
rect -159 495 -153 501
rect -147 495 -141 501
rect -135 495 -129 501
rect -123 495 -117 501
rect -111 495 -105 501
rect -99 495 -93 501
rect -87 495 -81 501
rect -75 495 -69 501
rect -63 495 -57 501
rect -51 495 -45 501
rect -39 495 -33 501
rect -27 495 -21 501
rect -15 495 -9 501
rect -3 495 3 501
rect 9 495 15 501
rect 21 495 27 501
rect 33 495 39 501
rect 45 495 51 501
rect 57 495 63 501
rect 69 495 75 501
rect 81 495 87 501
rect 93 495 99 501
rect 105 495 111 501
rect 117 495 123 501
rect 129 495 135 501
rect 141 495 147 501
rect 153 495 159 501
rect 165 495 171 501
rect 177 495 183 501
rect 189 495 195 501
rect 201 495 207 501
rect 213 495 219 501
rect 225 495 231 501
rect 237 495 243 501
rect 249 495 255 501
rect 261 495 264 501
rect -372 492 264 495
rect 276 597 288 603
rect 276 591 279 597
rect 285 591 288 597
rect 276 585 288 591
rect 276 579 279 585
rect 285 579 288 585
rect 276 573 288 579
rect 276 567 279 573
rect 285 567 288 573
rect 276 561 288 567
rect 276 555 279 561
rect 285 555 288 561
rect 276 549 288 555
rect 276 543 279 549
rect 285 543 288 549
rect 276 537 288 543
rect 276 531 279 537
rect 285 531 288 537
rect 276 525 288 531
rect 276 519 279 525
rect 285 519 288 525
rect 276 513 288 519
rect 276 507 279 513
rect 285 507 288 513
rect 276 501 288 507
rect 276 495 279 501
rect 285 495 288 501
rect -396 483 -393 489
rect -387 483 -384 489
rect -396 480 -384 483
rect 276 489 288 495
rect 276 483 279 489
rect 285 483 288 489
rect 276 480 288 483
rect -396 477 288 480
rect -396 471 -393 477
rect -387 471 -381 477
rect -375 471 -369 477
rect -363 471 -357 477
rect -351 471 -345 477
rect -339 471 -333 477
rect -327 471 -321 477
rect -315 471 -309 477
rect -303 471 -297 477
rect -291 471 -285 477
rect -279 471 -273 477
rect -267 471 -261 477
rect -255 471 -249 477
rect -243 471 -237 477
rect -231 471 -225 477
rect -219 471 -213 477
rect -207 471 -201 477
rect -195 471 -189 477
rect -183 471 -177 477
rect -171 471 -165 477
rect -159 471 -153 477
rect -147 471 -141 477
rect -135 471 -129 477
rect -123 471 -117 477
rect -111 471 -105 477
rect -99 471 -93 477
rect -87 471 -81 477
rect -75 471 -69 477
rect -63 471 -57 477
rect -51 471 -45 477
rect -39 471 -33 477
rect -27 471 -21 477
rect -15 471 -9 477
rect -3 471 3 477
rect 9 471 15 477
rect 21 471 27 477
rect 33 471 39 477
rect 45 471 51 477
rect 57 471 63 477
rect 69 471 75 477
rect 81 471 87 477
rect 93 471 99 477
rect 105 471 111 477
rect 117 471 123 477
rect 129 471 135 477
rect 141 471 147 477
rect 153 471 159 477
rect 165 471 171 477
rect 177 471 183 477
rect 189 471 195 477
rect 201 471 207 477
rect 213 471 219 477
rect 225 471 231 477
rect 237 471 243 477
rect 249 471 255 477
rect 261 471 267 477
rect 273 471 279 477
rect 285 471 288 477
rect -396 468 288 471
rect -396 465 -384 468
rect -396 459 -393 465
rect -387 459 -384 465
rect -396 453 -384 459
rect 276 465 288 468
rect 276 459 279 465
rect 285 459 288 465
rect -396 447 -393 453
rect -387 447 -384 453
rect -396 441 -384 447
rect -396 435 -393 441
rect -387 435 -384 441
rect -396 429 -384 435
rect -396 423 -393 429
rect -387 423 -384 429
rect -396 417 -384 423
rect -396 411 -393 417
rect -387 411 -384 417
rect -396 405 -384 411
rect -396 399 -393 405
rect -387 399 -384 405
rect -396 393 -384 399
rect -396 387 -393 393
rect -387 387 -384 393
rect -396 381 -384 387
rect -396 375 -393 381
rect -387 375 -384 381
rect -396 369 -384 375
rect -396 363 -393 369
rect -387 363 -384 369
rect -396 357 -384 363
rect -396 351 -393 357
rect -387 351 -384 357
rect -396 345 -384 351
rect -372 453 264 456
rect -372 447 -369 453
rect -363 447 -357 453
rect -351 447 -345 453
rect -339 447 -333 453
rect -327 447 -321 453
rect -315 447 -309 453
rect -303 447 -297 453
rect -291 447 -285 453
rect -279 447 -273 453
rect -267 447 -261 453
rect -255 447 -249 453
rect -243 447 -237 453
rect -231 447 -225 453
rect -219 447 -213 453
rect -207 447 -201 453
rect -195 447 -189 453
rect -183 447 -177 453
rect -171 447 -165 453
rect -159 447 -153 453
rect -147 447 -141 453
rect -135 447 -129 453
rect -123 447 -117 453
rect -111 447 -105 453
rect -99 447 -93 453
rect -87 447 -81 453
rect -75 447 -69 453
rect -63 447 -57 453
rect -51 447 -45 453
rect -39 447 -33 453
rect -27 447 -21 453
rect -15 447 -9 453
rect -3 447 3 453
rect 9 447 15 453
rect 21 447 27 453
rect 33 447 39 453
rect 45 447 51 453
rect 57 447 63 453
rect 69 447 75 453
rect 81 447 87 453
rect 93 447 99 453
rect 105 447 111 453
rect 117 447 123 453
rect 129 447 135 453
rect 141 447 147 453
rect 153 447 159 453
rect 165 447 171 453
rect 177 447 183 453
rect 189 447 195 453
rect 201 447 207 453
rect 213 447 219 453
rect 225 447 231 453
rect 237 447 243 453
rect 249 447 255 453
rect 261 447 264 453
rect -372 444 264 447
rect -372 441 -360 444
rect -372 435 -369 441
rect -363 435 -360 441
rect -372 429 -360 435
rect 252 441 264 444
rect 252 435 255 441
rect 261 435 264 441
rect -372 423 -369 429
rect -363 423 -360 429
rect -372 417 -360 423
rect -372 411 -369 417
rect -363 411 -360 417
rect -372 405 -360 411
rect -372 399 -369 405
rect -363 399 -360 405
rect -372 393 -360 399
rect -348 429 -336 432
rect -348 423 -345 429
rect -339 423 -336 429
rect -348 417 -336 423
rect -300 429 -288 432
rect -300 423 -297 429
rect -291 423 -288 429
rect -348 411 -345 417
rect -339 411 -336 417
rect -348 405 -336 411
rect -348 399 -345 405
rect -339 399 -336 405
rect -348 396 -336 399
rect -324 417 -312 420
rect -324 411 -321 417
rect -315 411 -312 417
rect -324 405 -312 411
rect -324 399 -321 405
rect -315 399 -312 405
rect -324 396 -312 399
rect -300 417 -288 423
rect -252 429 -240 432
rect -252 423 -249 429
rect -243 423 -240 429
rect -300 411 -297 417
rect -291 411 -288 417
rect -300 405 -288 411
rect -300 399 -297 405
rect -291 399 -288 405
rect -300 396 -288 399
rect -276 417 -264 420
rect -276 411 -273 417
rect -267 411 -264 417
rect -276 405 -264 411
rect -276 399 -273 405
rect -267 399 -264 405
rect -276 396 -264 399
rect -252 417 -240 423
rect -204 429 -192 432
rect -204 423 -201 429
rect -195 423 -192 429
rect -252 411 -249 417
rect -243 411 -240 417
rect -252 405 -240 411
rect -252 399 -249 405
rect -243 399 -240 405
rect -252 396 -240 399
rect -228 417 -216 420
rect -228 411 -225 417
rect -219 411 -216 417
rect -228 405 -216 411
rect -228 399 -225 405
rect -219 399 -216 405
rect -228 396 -216 399
rect -204 417 -192 423
rect -156 429 -144 432
rect -156 423 -153 429
rect -147 423 -144 429
rect -204 411 -201 417
rect -195 411 -192 417
rect -204 405 -192 411
rect -204 399 -201 405
rect -195 399 -192 405
rect -204 396 -192 399
rect -180 417 -168 420
rect -180 411 -177 417
rect -171 411 -168 417
rect -180 405 -168 411
rect -180 399 -177 405
rect -171 399 -168 405
rect -180 396 -168 399
rect -156 417 -144 423
rect -108 429 -96 432
rect -108 423 -105 429
rect -99 423 -96 429
rect -156 411 -153 417
rect -147 411 -144 417
rect -156 405 -144 411
rect -156 399 -153 405
rect -147 399 -144 405
rect -156 396 -144 399
rect -132 417 -120 420
rect -132 411 -129 417
rect -123 411 -120 417
rect -132 405 -120 411
rect -132 399 -129 405
rect -123 399 -120 405
rect -132 396 -120 399
rect -108 417 -96 423
rect -60 429 -48 432
rect -60 423 -57 429
rect -51 423 -48 429
rect -108 411 -105 417
rect -99 411 -96 417
rect -108 405 -96 411
rect -108 399 -105 405
rect -99 399 -96 405
rect -108 396 -96 399
rect -84 417 -72 420
rect -84 411 -81 417
rect -75 411 -72 417
rect -84 405 -72 411
rect -84 399 -81 405
rect -75 399 -72 405
rect -84 396 -72 399
rect -60 417 -48 423
rect -12 429 0 432
rect -12 423 -9 429
rect -3 423 0 429
rect -60 411 -57 417
rect -51 411 -48 417
rect -60 405 -48 411
rect -60 399 -57 405
rect -51 399 -48 405
rect -60 396 -48 399
rect -36 417 -24 420
rect -36 411 -33 417
rect -27 411 -24 417
rect -36 405 -24 411
rect -36 399 -33 405
rect -27 399 -24 405
rect -36 396 -24 399
rect -12 417 0 423
rect 36 429 48 432
rect 36 423 39 429
rect 45 423 48 429
rect -12 411 -9 417
rect -3 411 0 417
rect -12 405 0 411
rect -12 399 -9 405
rect -3 399 0 405
rect -12 396 0 399
rect 12 417 24 420
rect 12 411 15 417
rect 21 411 24 417
rect 12 405 24 411
rect 12 399 15 405
rect 21 399 24 405
rect 12 396 24 399
rect 36 417 48 423
rect 84 429 96 432
rect 84 423 87 429
rect 93 423 96 429
rect 36 411 39 417
rect 45 411 48 417
rect 36 405 48 411
rect 36 399 39 405
rect 45 399 48 405
rect 36 396 48 399
rect 60 417 72 420
rect 60 411 63 417
rect 69 411 72 417
rect 60 405 72 411
rect 60 399 63 405
rect 69 399 72 405
rect 60 396 72 399
rect 84 417 96 423
rect 132 429 144 432
rect 132 423 135 429
rect 141 423 144 429
rect 84 411 87 417
rect 93 411 96 417
rect 84 405 96 411
rect 84 399 87 405
rect 93 399 96 405
rect 84 396 96 399
rect 108 417 120 420
rect 108 411 111 417
rect 117 411 120 417
rect 108 405 120 411
rect 108 399 111 405
rect 117 399 120 405
rect 108 396 120 399
rect 132 417 144 423
rect 180 429 192 432
rect 180 423 183 429
rect 189 423 192 429
rect 132 411 135 417
rect 141 411 144 417
rect 132 405 144 411
rect 132 399 135 405
rect 141 399 144 405
rect 132 396 144 399
rect 156 417 168 420
rect 156 411 159 417
rect 165 411 168 417
rect 156 405 168 411
rect 156 399 159 405
rect 165 399 168 405
rect 156 396 168 399
rect 180 417 192 423
rect 228 429 240 432
rect 228 423 231 429
rect 237 423 240 429
rect 180 411 183 417
rect 189 411 192 417
rect 180 405 192 411
rect 180 399 183 405
rect 189 399 192 405
rect 180 396 192 399
rect 204 417 216 420
rect 204 411 207 417
rect 213 411 216 417
rect 204 405 216 411
rect 204 399 207 405
rect 213 399 216 405
rect 204 396 216 399
rect 228 417 240 423
rect 228 411 231 417
rect 237 411 240 417
rect 228 405 240 411
rect 228 399 231 405
rect 237 399 240 405
rect 228 396 240 399
rect 252 429 264 435
rect 252 423 255 429
rect 261 423 264 429
rect 252 417 264 423
rect 252 411 255 417
rect 261 411 264 417
rect 252 405 264 411
rect 252 399 255 405
rect 261 399 264 405
rect -372 387 -369 393
rect -363 387 -360 393
rect -372 381 -360 387
rect 252 393 264 399
rect 252 387 255 393
rect 261 387 264 393
rect -372 375 -369 381
rect -363 375 -360 381
rect -372 369 -360 375
rect -336 381 -300 384
rect -336 375 -333 381
rect -327 375 -321 381
rect -315 375 -309 381
rect -303 375 -300 381
rect -336 372 -300 375
rect -288 381 -252 384
rect -288 375 -285 381
rect -279 375 -273 381
rect -267 375 -261 381
rect -255 375 -252 381
rect -288 372 -252 375
rect -240 381 -204 384
rect -240 375 -237 381
rect -231 375 -225 381
rect -219 375 -213 381
rect -207 375 -204 381
rect -240 372 -204 375
rect -192 381 -156 384
rect -192 375 -189 381
rect -183 375 -177 381
rect -171 375 -165 381
rect -159 375 -156 381
rect -192 372 -156 375
rect -144 381 -108 384
rect -144 375 -141 381
rect -135 375 -129 381
rect -123 375 -117 381
rect -111 375 -108 381
rect -144 372 -108 375
rect -96 381 -60 384
rect -96 375 -93 381
rect -87 375 -81 381
rect -75 375 -69 381
rect -63 375 -60 381
rect -96 372 -60 375
rect -48 381 -12 384
rect -48 375 -45 381
rect -39 375 -33 381
rect -27 375 -21 381
rect -15 375 -12 381
rect -48 372 -12 375
rect 0 381 36 384
rect 0 375 3 381
rect 9 375 15 381
rect 21 375 27 381
rect 33 375 36 381
rect 0 372 36 375
rect 48 381 84 384
rect 48 375 51 381
rect 57 375 63 381
rect 69 375 75 381
rect 81 375 84 381
rect 48 372 84 375
rect 96 381 132 384
rect 96 375 99 381
rect 105 375 111 381
rect 117 375 123 381
rect 129 375 132 381
rect 96 372 132 375
rect 144 381 180 384
rect 144 375 147 381
rect 153 375 159 381
rect 165 375 171 381
rect 177 375 180 381
rect 144 372 180 375
rect 192 381 228 384
rect 192 375 195 381
rect 201 375 207 381
rect 213 375 219 381
rect 225 375 228 381
rect 192 372 228 375
rect 252 381 264 387
rect 252 375 255 381
rect 261 375 264 381
rect -372 363 -369 369
rect -363 363 -360 369
rect -372 360 -360 363
rect 252 369 264 375
rect 252 363 255 369
rect 261 363 264 369
rect 252 360 264 363
rect -372 357 264 360
rect -372 351 -369 357
rect -363 351 -357 357
rect -351 351 -345 357
rect -339 351 -333 357
rect -327 351 -321 357
rect -315 351 -309 357
rect -303 351 -297 357
rect -291 351 -285 357
rect -279 351 -273 357
rect -267 351 -261 357
rect -255 351 -249 357
rect -243 351 -237 357
rect -231 351 -225 357
rect -219 351 -213 357
rect -207 351 -201 357
rect -195 351 -189 357
rect -183 351 -177 357
rect -171 351 -165 357
rect -159 351 -153 357
rect -147 351 -141 357
rect -135 351 -129 357
rect -123 351 -117 357
rect -111 351 -105 357
rect -99 351 -93 357
rect -87 351 -81 357
rect -75 351 -69 357
rect -63 351 -57 357
rect -51 351 -45 357
rect -39 351 -33 357
rect -27 351 -21 357
rect -15 351 -9 357
rect -3 351 3 357
rect 9 351 15 357
rect 21 351 27 357
rect 33 351 39 357
rect 45 351 51 357
rect 57 351 63 357
rect 69 351 75 357
rect 81 351 87 357
rect 93 351 99 357
rect 105 351 111 357
rect 117 351 123 357
rect 129 351 135 357
rect 141 351 147 357
rect 153 351 159 357
rect 165 351 171 357
rect 177 351 183 357
rect 189 351 195 357
rect 201 351 207 357
rect 213 351 219 357
rect 225 351 231 357
rect 237 351 243 357
rect 249 351 255 357
rect 261 351 264 357
rect -372 348 264 351
rect 276 453 288 459
rect 276 447 279 453
rect 285 447 288 453
rect 276 441 288 447
rect 276 435 279 441
rect 285 435 288 441
rect 276 429 288 435
rect 276 423 279 429
rect 285 423 288 429
rect 276 417 288 423
rect 276 411 279 417
rect 285 411 288 417
rect 276 405 288 411
rect 276 399 279 405
rect 285 399 288 405
rect 276 393 288 399
rect 276 387 279 393
rect 285 387 288 393
rect 276 381 288 387
rect 276 375 279 381
rect 285 375 288 381
rect 276 369 288 375
rect 276 363 279 369
rect 285 363 288 369
rect 276 357 288 363
rect 276 351 279 357
rect 285 351 288 357
rect -396 339 -393 345
rect -387 339 -384 345
rect -396 336 -384 339
rect 276 345 288 351
rect 276 339 279 345
rect 285 339 288 345
rect 276 336 288 339
rect -396 333 288 336
rect -396 327 -393 333
rect -387 327 -381 333
rect -375 327 -369 333
rect -363 327 -357 333
rect -351 327 -345 333
rect -339 327 -333 333
rect -327 327 -321 333
rect -315 327 -309 333
rect -303 327 -297 333
rect -291 327 -285 333
rect -279 327 -273 333
rect -267 327 -261 333
rect -255 327 -249 333
rect -243 327 -237 333
rect -231 327 -225 333
rect -219 327 -213 333
rect -207 327 -201 333
rect -195 327 -189 333
rect -183 327 -177 333
rect -171 327 -165 333
rect -159 327 -153 333
rect -147 327 -141 333
rect -135 327 -129 333
rect -123 327 -117 333
rect -111 327 -105 333
rect -99 327 -93 333
rect -87 327 -81 333
rect -75 327 -69 333
rect -63 327 -57 333
rect -51 327 -45 333
rect -39 327 -33 333
rect -27 327 -21 333
rect -15 327 -9 333
rect -3 327 3 333
rect 9 327 15 333
rect 21 327 27 333
rect 33 327 39 333
rect 45 327 51 333
rect 57 327 63 333
rect 69 327 75 333
rect 81 327 87 333
rect 93 327 99 333
rect 105 327 111 333
rect 117 327 123 333
rect 129 327 135 333
rect 141 327 147 333
rect 153 327 159 333
rect 165 327 171 333
rect 177 327 183 333
rect 189 327 195 333
rect 201 327 207 333
rect 213 327 219 333
rect 225 327 231 333
rect 237 327 243 333
rect 249 327 255 333
rect 261 327 267 333
rect 273 327 279 333
rect 285 327 288 333
rect -396 324 288 327
rect -396 321 -384 324
rect -396 315 -393 321
rect -387 315 -384 321
rect -396 309 -384 315
rect -396 303 -393 309
rect -387 303 -384 309
rect -396 297 -384 303
rect -396 291 -393 297
rect -387 291 -384 297
rect -396 285 -384 291
rect -396 279 -393 285
rect -387 279 -384 285
rect -396 273 -384 279
rect -396 267 -393 273
rect -387 267 -384 273
rect -396 261 -384 267
rect -396 255 -393 261
rect -387 255 -384 261
rect -396 249 -384 255
rect -396 243 -393 249
rect -387 243 -384 249
rect -396 237 -384 243
rect -396 231 -393 237
rect -387 231 -384 237
rect -396 225 -384 231
rect -396 219 -393 225
rect -387 219 -384 225
rect -396 213 -384 219
rect -396 207 -393 213
rect -387 207 -384 213
rect -396 201 -384 207
rect -396 195 -393 201
rect -387 195 -384 201
rect -396 189 -384 195
rect -396 183 -393 189
rect -387 183 -384 189
rect -396 177 -384 183
rect -396 171 -393 177
rect -387 171 -384 177
rect -396 165 -384 171
rect -396 159 -393 165
rect -387 159 -384 165
rect -396 153 -384 159
rect -396 147 -393 153
rect -387 147 -384 153
rect -396 141 -384 147
rect -396 135 -393 141
rect -387 135 -384 141
rect -396 129 -384 135
rect -396 123 -393 129
rect -387 123 -384 129
rect -396 117 -384 123
rect -396 111 -393 117
rect -387 111 -384 117
rect -396 105 -384 111
rect -396 99 -393 105
rect -387 99 -384 105
rect -396 96 -384 99
rect 276 321 288 324
rect 276 315 279 321
rect 285 315 288 321
rect 276 309 288 315
rect 276 303 279 309
rect 285 303 288 309
rect 276 297 288 303
rect 276 291 279 297
rect 285 291 288 297
rect 276 285 288 291
rect 276 279 279 285
rect 285 279 288 285
rect 276 273 288 279
rect 276 267 279 273
rect 285 267 288 273
rect 276 261 288 267
rect 276 255 279 261
rect 285 255 288 261
rect 276 249 288 255
rect 276 243 279 249
rect 285 243 288 249
rect 276 237 288 243
rect 276 231 279 237
rect 285 231 288 237
rect 276 225 288 231
rect 276 219 279 225
rect 285 219 288 225
rect 276 213 288 219
rect 276 207 279 213
rect 285 207 288 213
rect 276 201 288 207
rect 276 195 279 201
rect 285 195 288 201
rect 276 189 288 195
rect 276 183 279 189
rect 285 183 288 189
rect 276 177 288 183
rect 276 171 279 177
rect 285 171 288 177
rect 276 165 288 171
rect 276 159 279 165
rect 285 159 288 165
rect 276 153 288 159
rect 276 147 279 153
rect 285 147 288 153
rect 276 141 288 147
rect 276 135 279 141
rect 285 135 288 141
rect 276 129 288 135
rect 276 123 279 129
rect 285 123 288 129
rect 276 117 288 123
rect 276 111 279 117
rect 285 111 288 117
rect 276 105 288 111
rect 276 99 279 105
rect 285 99 288 105
rect 276 96 288 99
rect -396 93 288 96
rect -396 87 -393 93
rect -387 87 -381 93
rect -375 87 -369 93
rect -363 87 -357 93
rect -351 87 -345 93
rect -339 87 -333 93
rect -327 87 -321 93
rect -315 87 -309 93
rect -303 87 -297 93
rect -291 87 -285 93
rect -279 87 -273 93
rect -267 87 -261 93
rect -255 87 -249 93
rect -243 87 -237 93
rect -231 87 -225 93
rect -219 87 -213 93
rect -207 87 -201 93
rect -195 87 -189 93
rect -183 87 -177 93
rect -171 87 -165 93
rect -159 87 -153 93
rect -147 87 -141 93
rect -135 87 -129 93
rect -123 87 -117 93
rect -111 87 -105 93
rect -99 87 -93 93
rect -87 87 -81 93
rect -75 87 -69 93
rect -63 87 -57 93
rect -51 87 -45 93
rect -39 87 -33 93
rect -27 87 -21 93
rect -15 87 -9 93
rect -3 87 3 93
rect 9 87 15 93
rect 21 87 27 93
rect 33 87 39 93
rect 45 87 51 93
rect 57 87 63 93
rect 69 87 75 93
rect 81 87 87 93
rect 93 87 99 93
rect 105 87 111 93
rect 117 87 123 93
rect 129 87 135 93
rect 141 87 147 93
rect 153 87 159 93
rect 165 87 171 93
rect 177 87 183 93
rect 189 87 195 93
rect 201 87 207 93
rect 213 87 219 93
rect 225 87 231 93
rect 237 87 243 93
rect 249 87 255 93
rect 261 87 267 93
rect 273 87 279 93
rect 285 87 288 93
rect -396 84 288 87
rect -396 81 -384 84
rect -396 75 -393 81
rect -387 75 -384 81
rect -396 69 -384 75
rect 276 81 288 84
rect 276 75 279 81
rect 285 75 288 81
rect -396 63 -393 69
rect -387 63 -384 69
rect -396 57 -384 63
rect -336 69 -300 72
rect -336 63 -333 69
rect -327 63 -321 69
rect -315 63 -309 69
rect -303 63 -300 69
rect -336 60 -300 63
rect -288 69 -252 72
rect -288 63 -285 69
rect -279 63 -273 69
rect -267 63 -261 69
rect -255 63 -252 69
rect -288 60 -252 63
rect -240 69 -204 72
rect -240 63 -237 69
rect -231 63 -225 69
rect -219 63 -213 69
rect -207 63 -204 69
rect -240 60 -204 63
rect -192 69 -156 72
rect -192 63 -189 69
rect -183 63 -177 69
rect -171 63 -165 69
rect -159 63 -156 69
rect -192 60 -156 63
rect -144 69 -108 72
rect -144 63 -141 69
rect -135 63 -129 69
rect -123 63 -117 69
rect -111 63 -108 69
rect -144 60 -108 63
rect -96 69 -60 72
rect -96 63 -93 69
rect -87 63 -81 69
rect -75 63 -69 69
rect -63 63 -60 69
rect -96 60 -60 63
rect -48 69 -12 72
rect -48 63 -45 69
rect -39 63 -33 69
rect -27 63 -21 69
rect -15 63 -12 69
rect -48 60 -12 63
rect 0 69 36 72
rect 0 63 3 69
rect 9 63 15 69
rect 21 63 27 69
rect 33 63 36 69
rect 0 60 36 63
rect 48 69 84 72
rect 48 63 51 69
rect 57 63 63 69
rect 69 63 75 69
rect 81 63 84 69
rect 48 60 84 63
rect 96 69 132 72
rect 96 63 99 69
rect 105 63 111 69
rect 117 63 123 69
rect 129 63 132 69
rect 96 60 132 63
rect 144 69 180 72
rect 144 63 147 69
rect 153 63 159 69
rect 165 63 171 69
rect 177 63 180 69
rect 144 60 180 63
rect 192 69 228 72
rect 192 63 195 69
rect 201 63 207 69
rect 213 63 219 69
rect 225 63 228 69
rect 192 60 228 63
rect 276 69 288 75
rect 276 63 279 69
rect 285 63 288 69
rect -396 51 -393 57
rect -387 51 -384 57
rect -396 45 -384 51
rect -396 39 -393 45
rect -387 39 -384 45
rect -396 33 -384 39
rect -396 27 -393 33
rect -387 27 -384 33
rect -396 21 -384 27
rect -396 15 -393 21
rect -387 15 -384 21
rect -396 9 -384 15
rect -348 45 -336 48
rect -348 39 -345 45
rect -339 39 -336 45
rect -348 33 -336 39
rect -348 27 -345 33
rect -339 27 -336 33
rect -348 21 -336 27
rect -348 15 -345 21
rect -339 15 -336 21
rect -348 12 -336 15
rect -324 45 -312 60
rect 276 57 288 63
rect 276 51 279 57
rect 285 51 288 57
rect -324 39 -321 45
rect -315 39 -312 45
rect -324 33 -312 39
rect -324 27 -321 33
rect -315 27 -312 33
rect -324 21 -312 27
rect -324 15 -321 21
rect -315 15 -312 21
rect -324 12 -312 15
rect -300 45 -288 48
rect -300 39 -297 45
rect -291 39 -288 45
rect -300 33 -288 39
rect -300 27 -297 33
rect -291 27 -288 33
rect -300 21 -288 27
rect -300 15 -297 21
rect -291 15 -288 21
rect -300 12 -288 15
rect -276 45 -264 48
rect -276 39 -273 45
rect -267 39 -264 45
rect -276 33 -264 39
rect -276 27 -273 33
rect -267 27 -264 33
rect -276 21 -264 27
rect -276 15 -273 21
rect -267 15 -264 21
rect -276 12 -264 15
rect -252 45 -240 48
rect -252 39 -249 45
rect -243 39 -240 45
rect -252 33 -240 39
rect -252 27 -249 33
rect -243 27 -240 33
rect -252 21 -240 27
rect -252 15 -249 21
rect -243 15 -240 21
rect -252 12 -240 15
rect -228 45 -216 48
rect -228 39 -225 45
rect -219 39 -216 45
rect -228 33 -216 39
rect -228 27 -225 33
rect -219 27 -216 33
rect -228 21 -216 27
rect -228 15 -225 21
rect -219 15 -216 21
rect -228 12 -216 15
rect -204 45 -192 48
rect -204 39 -201 45
rect -195 39 -192 45
rect -204 33 -192 39
rect -204 27 -201 33
rect -195 27 -192 33
rect -204 21 -192 27
rect -204 15 -201 21
rect -195 15 -192 21
rect -204 12 -192 15
rect -180 45 -168 48
rect -180 39 -177 45
rect -171 39 -168 45
rect -180 33 -168 39
rect -180 27 -177 33
rect -171 27 -168 33
rect -180 21 -168 27
rect -180 15 -177 21
rect -171 15 -168 21
rect -180 12 -168 15
rect -156 45 -144 48
rect -156 39 -153 45
rect -147 39 -144 45
rect -156 33 -144 39
rect -156 27 -153 33
rect -147 27 -144 33
rect -156 21 -144 27
rect -156 15 -153 21
rect -147 15 -144 21
rect -156 12 -144 15
rect -132 45 -120 48
rect -132 39 -129 45
rect -123 39 -120 45
rect -132 33 -120 39
rect -132 27 -129 33
rect -123 27 -120 33
rect -132 21 -120 27
rect -132 15 -129 21
rect -123 15 -120 21
rect -132 12 -120 15
rect -108 45 -96 48
rect -108 39 -105 45
rect -99 39 -96 45
rect -108 33 -96 39
rect -108 27 -105 33
rect -99 27 -96 33
rect -108 21 -96 27
rect -108 15 -105 21
rect -99 15 -96 21
rect -108 12 -96 15
rect -60 45 -48 48
rect -60 39 -57 45
rect -51 39 -48 45
rect -60 33 -48 39
rect -60 27 -57 33
rect -51 27 -48 33
rect -60 21 -48 27
rect -60 15 -57 21
rect -51 15 -48 21
rect -60 12 -48 15
rect -12 45 0 48
rect -12 39 -9 45
rect -3 39 0 45
rect -12 33 0 39
rect -12 27 -9 33
rect -3 27 0 33
rect -12 21 0 27
rect -12 15 -9 21
rect -3 15 0 21
rect -12 12 0 15
rect 36 45 48 48
rect 36 39 39 45
rect 45 39 48 45
rect 36 33 48 39
rect 36 27 39 33
rect 45 27 48 33
rect 36 21 48 27
rect 36 15 39 21
rect 45 15 48 21
rect 36 12 48 15
rect 84 45 96 48
rect 84 39 87 45
rect 93 39 96 45
rect 84 33 96 39
rect 84 27 87 33
rect 93 27 96 33
rect 84 21 96 27
rect 84 15 87 21
rect 93 15 96 21
rect 84 12 96 15
rect 132 45 144 48
rect 132 39 135 45
rect 141 39 144 45
rect 132 33 144 39
rect 132 27 135 33
rect 141 27 144 33
rect 132 21 144 27
rect 132 15 135 21
rect 141 15 144 21
rect 132 12 144 15
rect 180 45 192 48
rect 180 39 183 45
rect 189 39 192 45
rect 180 33 192 39
rect 180 27 183 33
rect 189 27 192 33
rect 180 21 192 27
rect 180 15 183 21
rect 189 15 192 21
rect 180 12 192 15
rect 204 45 216 48
rect 204 39 207 45
rect 213 39 216 45
rect 204 33 216 39
rect 204 27 207 33
rect 213 27 216 33
rect 204 21 216 27
rect 204 15 207 21
rect 213 15 216 21
rect 204 12 216 15
rect 228 45 240 48
rect 228 39 231 45
rect 237 39 240 45
rect 228 33 240 39
rect 228 27 231 33
rect 237 27 240 33
rect 228 21 240 27
rect 228 15 231 21
rect 237 15 240 21
rect 228 12 240 15
rect 276 45 288 51
rect 276 39 279 45
rect 285 39 288 45
rect 276 33 288 39
rect 276 27 279 33
rect 285 27 288 33
rect 276 21 288 27
rect 276 15 279 21
rect 285 15 288 21
rect -396 3 -393 9
rect -387 3 -384 9
rect -396 0 -384 3
rect 276 9 288 15
rect 276 3 279 9
rect 285 3 288 9
rect 276 0 288 3
rect -396 -3 288 0
rect -396 -9 -393 -3
rect -387 -9 -381 -3
rect -375 -9 -369 -3
rect -363 -9 -357 -3
rect -351 -9 -345 -3
rect -339 -9 -333 -3
rect -327 -9 -321 -3
rect -315 -9 -309 -3
rect -303 -9 -297 -3
rect -291 -9 -285 -3
rect -279 -9 -273 -3
rect -267 -9 -261 -3
rect -255 -9 -249 -3
rect -243 -9 -237 -3
rect -231 -9 -225 -3
rect -219 -9 -213 -3
rect -207 -9 -201 -3
rect -195 -9 -189 -3
rect -183 -9 -177 -3
rect -171 -9 -165 -3
rect -159 -9 -153 -3
rect -147 -9 -141 -3
rect -135 -9 -129 -3
rect -123 -9 -117 -3
rect -111 -9 -105 -3
rect -99 -9 -93 -3
rect -87 -9 -81 -3
rect -75 -9 -69 -3
rect -63 -9 -57 -3
rect -51 -9 -45 -3
rect -39 -9 -33 -3
rect -27 -9 -21 -3
rect -15 -9 -9 -3
rect -3 -9 3 -3
rect 9 -9 15 -3
rect 21 -9 27 -3
rect 33 -9 39 -3
rect 45 -9 51 -3
rect 57 -9 63 -3
rect 69 -9 75 -3
rect 81 -9 87 -3
rect 93 -9 99 -3
rect 105 -9 111 -3
rect 117 -9 123 -3
rect 129 -9 135 -3
rect 141 -9 147 -3
rect 153 -9 159 -3
rect 165 -9 171 -3
rect 177 -9 183 -3
rect 189 -9 195 -3
rect 201 -9 207 -3
rect 213 -9 219 -3
rect 225 -9 231 -3
rect 237 -9 243 -3
rect 249 -9 255 -3
rect 261 -9 267 -3
rect 273 -9 279 -3
rect 285 -9 288 -3
rect -396 -12 288 -9
<< via1 >>
rect -321 567 -315 573
rect -273 567 -267 573
rect -225 567 -219 573
rect -177 567 -171 573
rect -129 567 -123 573
rect -81 567 -75 573
rect -33 567 -27 573
rect 15 567 21 573
rect 63 567 69 573
rect 111 567 117 573
rect 159 567 165 573
rect 207 567 213 573
rect -345 543 -339 549
rect -345 531 -339 537
rect -345 519 -339 525
rect -321 543 -315 549
rect -321 531 -315 537
rect -321 519 -315 525
rect -297 543 -291 549
rect -297 531 -291 537
rect -297 519 -291 525
rect -273 543 -267 549
rect -273 531 -267 537
rect -273 519 -267 525
rect -249 543 -243 549
rect -249 531 -243 537
rect -249 519 -243 525
rect -225 543 -219 549
rect -225 531 -219 537
rect -225 519 -219 525
rect -201 543 -195 549
rect -201 531 -195 537
rect -201 519 -195 525
rect -177 543 -171 549
rect -177 531 -171 537
rect -177 519 -171 525
rect -153 543 -147 549
rect -153 531 -147 537
rect -153 519 -147 525
rect -129 543 -123 549
rect -129 531 -123 537
rect -129 519 -123 525
rect -105 543 -99 549
rect -105 531 -99 537
rect -105 519 -99 525
rect -81 543 -75 549
rect -81 531 -75 537
rect -81 519 -75 525
rect -57 543 -51 549
rect -57 531 -51 537
rect -57 519 -51 525
rect -33 543 -27 549
rect -33 531 -27 537
rect -33 519 -27 525
rect -9 543 -3 549
rect -9 531 -3 537
rect -9 519 -3 525
rect 15 543 21 549
rect 15 531 21 537
rect 15 519 21 525
rect 39 543 45 549
rect 39 531 45 537
rect 39 519 45 525
rect 63 543 69 549
rect 63 531 69 537
rect 63 519 69 525
rect 87 543 93 549
rect 87 531 93 537
rect 87 519 93 525
rect 111 543 117 549
rect 111 531 117 537
rect 111 519 117 525
rect 135 543 141 549
rect 135 531 141 537
rect 135 519 141 525
rect 159 543 165 549
rect 159 531 165 537
rect 159 519 165 525
rect 183 543 189 549
rect 183 531 189 537
rect 183 519 189 525
rect 207 543 213 549
rect 207 531 213 537
rect 207 519 213 525
rect 231 543 237 549
rect 231 531 237 537
rect 231 519 237 525
rect -225 447 -219 453
rect -177 447 -171 453
rect -345 423 -339 429
rect -297 423 -291 429
rect -345 411 -339 417
rect -345 399 -339 405
rect -321 399 -315 405
rect -249 423 -243 429
rect -201 423 -195 429
rect -225 399 -219 405
rect -153 423 -147 429
rect -177 399 -171 405
rect -105 423 -99 429
rect -153 411 -147 417
rect -153 399 -147 405
rect -57 423 -51 429
rect -105 411 -99 417
rect -105 399 -99 405
rect -81 399 -75 405
rect -9 423 -3 429
rect -33 399 -27 405
rect 39 423 45 429
rect -9 411 -3 417
rect -9 399 -3 405
rect 15 399 21 405
rect 87 423 93 429
rect 63 399 69 405
rect 135 423 141 429
rect 87 411 93 417
rect 87 399 93 405
rect 183 423 189 429
rect 135 411 141 417
rect 135 399 141 405
rect 231 423 237 429
rect 183 411 189 417
rect 183 399 189 405
rect 231 411 237 417
rect 231 399 237 405
rect -321 375 -315 381
rect -273 375 -267 381
rect -225 375 -219 381
rect -177 375 -171 381
rect -129 375 -123 381
rect -81 375 -75 381
rect -33 375 -27 381
rect 15 375 21 381
rect 63 375 69 381
rect 111 375 117 381
rect 159 375 165 381
rect 207 375 213 381
rect -345 327 -339 333
rect -297 327 -291 333
rect -153 327 -147 333
rect -105 327 -99 333
rect -9 327 -3 333
rect 87 327 93 333
rect 183 327 189 333
rect 231 327 237 333
rect -273 63 -267 69
rect -225 63 -219 69
rect -177 63 -171 69
rect -129 63 -123 69
rect -81 63 -75 69
rect -33 63 -27 69
rect 15 63 21 69
rect 63 63 69 69
rect 111 63 117 69
rect 159 63 165 69
rect 207 63 213 69
rect -345 39 -339 45
rect -345 27 -339 33
rect -345 15 -339 21
rect -321 39 -315 45
rect -321 27 -315 33
rect -321 15 -315 21
rect -297 39 -291 45
rect -297 27 -291 33
rect -297 15 -291 21
rect -273 39 -267 45
rect -273 27 -267 33
rect -273 15 -267 21
rect -249 15 -243 21
rect -201 39 -195 45
rect -201 27 -195 33
rect -201 15 -195 21
rect -153 39 -147 45
rect -153 27 -147 33
rect -153 15 -147 21
rect -105 39 -99 45
rect -105 27 -99 33
rect -105 15 -99 21
rect -57 39 -51 45
rect -57 27 -51 33
rect -57 15 -51 21
rect -9 39 -3 45
rect -9 27 -3 33
rect -9 15 -3 21
rect 39 39 45 45
rect 39 27 45 33
rect 39 15 45 21
rect 87 39 93 45
rect 87 27 93 33
rect 87 15 93 21
rect 135 39 141 45
rect 135 27 141 33
rect 135 15 141 21
rect 183 39 189 45
rect 183 27 189 33
rect 183 15 189 21
rect 231 39 237 45
rect 231 27 237 33
rect 231 15 237 21
rect -345 -9 -339 -3
rect -297 -9 -291 -3
rect -249 -9 -243 -3
rect -153 -9 -147 -3
rect -105 -9 -99 -3
rect -9 -9 -3 -3
rect 87 -9 93 -3
rect 183 -9 189 -3
rect 231 -9 237 -3
<< metal2 >>
rect -348 549 -336 600
rect -324 573 -312 576
rect -324 567 -321 573
rect -315 567 -312 573
rect -324 564 -312 567
rect -276 573 -264 576
rect -276 567 -273 573
rect -267 567 -264 573
rect -276 564 -264 567
rect -228 573 -216 576
rect -228 567 -225 573
rect -219 567 -216 573
rect -228 564 -216 567
rect -180 573 -168 576
rect -180 567 -177 573
rect -171 567 -168 573
rect -180 564 -168 567
rect -132 573 -120 576
rect -132 567 -129 573
rect -123 567 -120 573
rect -132 564 -120 567
rect -84 573 -72 576
rect -84 567 -81 573
rect -75 567 -72 573
rect -84 564 -72 567
rect -36 573 -24 576
rect -36 567 -33 573
rect -27 567 -24 573
rect -36 564 -24 567
rect 12 573 24 576
rect 12 567 15 573
rect 21 567 24 573
rect 12 564 24 567
rect 60 573 72 576
rect 60 567 63 573
rect 69 567 72 573
rect 60 564 72 567
rect 108 573 120 576
rect 108 567 111 573
rect 117 567 120 573
rect 108 564 120 567
rect 156 573 168 576
rect 156 567 159 573
rect 165 567 168 573
rect 156 564 168 567
rect 204 573 216 576
rect 204 567 207 573
rect 213 567 216 573
rect 204 564 216 567
rect -348 543 -345 549
rect -339 543 -336 549
rect -348 537 -336 543
rect -348 531 -345 537
rect -339 531 -336 537
rect -348 525 -336 531
rect -348 519 -345 525
rect -339 519 -336 525
rect -348 501 -336 519
rect -348 495 -345 501
rect -339 495 -336 501
rect -348 492 -336 495
rect -324 549 -312 552
rect -324 543 -321 549
rect -315 543 -312 549
rect -324 537 -312 543
rect -324 531 -321 537
rect -315 531 -312 537
rect -324 525 -312 531
rect -324 519 -321 525
rect -315 519 -312 525
rect -324 477 -312 519
rect -300 549 -288 552
rect -300 543 -297 549
rect -291 543 -288 549
rect -300 537 -288 543
rect -300 531 -297 537
rect -291 531 -288 537
rect -300 525 -288 531
rect -300 519 -297 525
rect -291 519 -288 525
rect -300 516 -288 519
rect -276 549 -264 552
rect -276 543 -273 549
rect -267 543 -264 549
rect -276 537 -264 543
rect -276 531 -273 537
rect -267 531 -264 537
rect -276 525 -264 531
rect -276 519 -273 525
rect -267 519 -264 525
rect -324 471 -321 477
rect -315 471 -312 477
rect -324 432 -312 471
rect -276 477 -264 519
rect -252 549 -240 552
rect -252 543 -249 549
rect -243 543 -240 549
rect -252 537 -240 543
rect -252 531 -249 537
rect -243 531 -240 537
rect -252 525 -240 531
rect -252 519 -249 525
rect -243 519 -240 525
rect -252 516 -240 519
rect -228 549 -216 552
rect -228 543 -225 549
rect -219 543 -216 549
rect -228 537 -216 543
rect -228 531 -225 537
rect -219 531 -216 537
rect -228 525 -216 531
rect -228 519 -225 525
rect -219 519 -216 525
rect -276 471 -273 477
rect -267 471 -264 477
rect -276 432 -264 471
rect -228 453 -216 519
rect -204 549 -192 552
rect -204 543 -201 549
rect -195 543 -192 549
rect -204 537 -192 543
rect -204 531 -201 537
rect -195 531 -192 537
rect -204 525 -192 531
rect -204 519 -201 525
rect -195 519 -192 525
rect -204 516 -192 519
rect -180 549 -168 552
rect -180 543 -177 549
rect -171 543 -168 549
rect -180 537 -168 543
rect -180 531 -177 537
rect -171 531 -168 537
rect -180 525 -168 531
rect -180 519 -177 525
rect -171 519 -168 525
rect -228 447 -225 453
rect -219 447 -216 453
rect -228 432 -216 447
rect -180 453 -168 519
rect -156 549 -144 552
rect -156 543 -153 549
rect -147 543 -144 549
rect -156 537 -144 543
rect -156 531 -153 537
rect -147 531 -144 537
rect -156 525 -144 531
rect -156 519 -153 525
rect -147 519 -144 525
rect -156 516 -144 519
rect -132 549 -120 552
rect -132 543 -129 549
rect -123 543 -120 549
rect -132 537 -120 543
rect -132 531 -129 537
rect -123 531 -120 537
rect -132 525 -120 531
rect -132 519 -129 525
rect -123 519 -120 525
rect -180 447 -177 453
rect -171 447 -168 453
rect -180 432 -168 447
rect -132 477 -120 519
rect -108 549 -96 552
rect -108 543 -105 549
rect -99 543 -96 549
rect -108 537 -96 543
rect -108 531 -105 537
rect -99 531 -96 537
rect -108 525 -96 531
rect -108 519 -105 525
rect -99 519 -96 525
rect -108 516 -96 519
rect -84 549 -72 552
rect -84 543 -81 549
rect -75 543 -72 549
rect -84 537 -72 543
rect -84 531 -81 537
rect -75 531 -72 537
rect -84 525 -72 531
rect -84 519 -81 525
rect -75 519 -72 525
rect -132 471 -129 477
rect -123 471 -120 477
rect -132 432 -120 471
rect -84 477 -72 519
rect -60 549 -48 552
rect -60 543 -57 549
rect -51 543 -48 549
rect -60 537 -48 543
rect -60 531 -57 537
rect -51 531 -48 537
rect -60 525 -48 531
rect -60 519 -57 525
rect -51 519 -48 525
rect -60 516 -48 519
rect -36 549 -24 552
rect -36 543 -33 549
rect -27 543 -24 549
rect -36 537 -24 543
rect -36 531 -33 537
rect -27 531 -24 537
rect -36 525 -24 531
rect -36 519 -33 525
rect -27 519 -24 525
rect -84 471 -81 477
rect -75 471 -72 477
rect -84 432 -72 471
rect -36 477 -24 519
rect -12 549 0 552
rect -12 543 -9 549
rect -3 543 0 549
rect -12 537 0 543
rect -12 531 -9 537
rect -3 531 0 537
rect -12 525 0 531
rect -12 519 -9 525
rect -3 519 0 525
rect -12 516 0 519
rect 12 549 24 552
rect 12 543 15 549
rect 21 543 24 549
rect 12 537 24 543
rect 12 531 15 537
rect 21 531 24 537
rect 12 525 24 531
rect 12 519 15 525
rect 21 519 24 525
rect -36 471 -33 477
rect -27 471 -24 477
rect -36 432 -24 471
rect 12 477 24 519
rect 36 549 48 552
rect 36 543 39 549
rect 45 543 48 549
rect 36 537 48 543
rect 36 531 39 537
rect 45 531 48 537
rect 36 525 48 531
rect 36 519 39 525
rect 45 519 48 525
rect 36 516 48 519
rect 60 549 72 552
rect 60 543 63 549
rect 69 543 72 549
rect 60 537 72 543
rect 60 531 63 537
rect 69 531 72 537
rect 60 525 72 531
rect 60 519 63 525
rect 69 519 72 525
rect 12 471 15 477
rect 21 471 24 477
rect 12 432 24 471
rect 60 477 72 519
rect 84 549 96 552
rect 84 543 87 549
rect 93 543 96 549
rect 84 537 96 543
rect 84 531 87 537
rect 93 531 96 537
rect 84 525 96 531
rect 84 519 87 525
rect 93 519 96 525
rect 84 516 96 519
rect 108 549 120 552
rect 108 543 111 549
rect 117 543 120 549
rect 108 537 120 543
rect 108 531 111 537
rect 117 531 120 537
rect 108 525 120 531
rect 108 519 111 525
rect 117 519 120 525
rect 60 471 63 477
rect 69 471 72 477
rect 60 432 72 471
rect 108 477 120 519
rect 132 549 144 552
rect 132 543 135 549
rect 141 543 144 549
rect 132 537 144 543
rect 132 531 135 537
rect 141 531 144 537
rect 132 525 144 531
rect 132 519 135 525
rect 141 519 144 525
rect 132 516 144 519
rect 156 549 168 552
rect 156 543 159 549
rect 165 543 168 549
rect 156 537 168 543
rect 156 531 159 537
rect 165 531 168 537
rect 156 525 168 531
rect 156 519 159 525
rect 165 519 168 525
rect 108 471 111 477
rect 117 471 120 477
rect 108 432 120 471
rect 156 477 168 519
rect 180 549 192 552
rect 180 543 183 549
rect 189 543 192 549
rect 180 537 192 543
rect 180 531 183 537
rect 189 531 192 537
rect 180 525 192 531
rect 180 519 183 525
rect 189 519 192 525
rect 180 516 192 519
rect 204 549 216 552
rect 204 543 207 549
rect 213 543 216 549
rect 204 537 216 543
rect 204 531 207 537
rect 213 531 216 537
rect 204 525 216 531
rect 204 519 207 525
rect 213 519 216 525
rect 156 471 159 477
rect 165 471 168 477
rect 156 432 168 471
rect 204 477 216 519
rect 228 549 240 552
rect 228 543 231 549
rect 237 543 240 549
rect 228 537 240 543
rect 228 531 231 537
rect 237 531 240 537
rect 228 525 240 531
rect 228 519 231 525
rect 237 519 240 525
rect 228 516 240 519
rect 204 471 207 477
rect 213 471 216 477
rect 204 432 216 471
rect -348 429 -264 432
rect -348 423 -345 429
rect -339 423 -297 429
rect -291 423 -264 429
rect -348 420 -264 423
rect -252 429 -144 432
rect -252 423 -249 429
rect -243 423 -201 429
rect -195 423 -153 429
rect -147 423 -144 429
rect -252 420 -144 423
rect -132 429 252 432
rect -132 423 -105 429
rect -99 423 -57 429
rect -51 423 -9 429
rect -3 423 39 429
rect 45 423 87 429
rect 93 423 135 429
rect 141 423 183 429
rect 189 423 231 429
rect 237 423 252 429
rect -132 420 252 423
rect -348 417 -336 420
rect -348 411 -345 417
rect -339 411 -336 417
rect -348 405 -336 411
rect -348 399 -345 405
rect -339 399 -336 405
rect -348 396 -336 399
rect -324 405 -264 408
rect -324 399 -321 405
rect -315 399 -264 405
rect -324 396 -264 399
rect -252 396 -240 420
rect -156 417 -144 420
rect -156 411 -153 417
rect -147 411 -144 417
rect -228 405 -168 408
rect -228 399 -225 405
rect -219 399 -177 405
rect -171 399 -168 405
rect -228 396 -168 399
rect -156 405 -144 411
rect -156 399 -153 405
rect -147 399 -144 405
rect -156 396 -144 399
rect -108 417 -96 420
rect -108 411 -105 417
rect -99 411 -96 417
rect -108 405 -96 411
rect -12 417 0 420
rect -12 411 -9 417
rect -3 411 0 417
rect -108 399 -105 405
rect -99 399 -96 405
rect -108 396 -96 399
rect -84 405 -24 408
rect -84 399 -81 405
rect -75 399 -33 405
rect -27 399 -24 405
rect -84 396 -24 399
rect -12 405 0 411
rect 84 417 96 420
rect 84 411 87 417
rect 93 411 96 417
rect -12 399 -9 405
rect -3 399 0 405
rect -12 396 0 399
rect 12 405 72 408
rect 12 399 15 405
rect 21 399 63 405
rect 69 399 72 405
rect 12 396 72 399
rect 84 405 96 411
rect 84 399 87 405
rect 93 399 96 405
rect 84 396 96 399
rect 132 417 144 420
rect 132 411 135 417
rect 141 411 144 417
rect 132 405 144 411
rect 132 399 135 405
rect 141 399 144 405
rect 132 396 144 399
rect 180 417 204 420
rect 180 411 183 417
rect 189 411 204 417
rect 180 405 204 411
rect 180 399 183 405
rect 189 399 204 405
rect 180 396 204 399
rect 228 417 252 420
rect 228 411 231 417
rect 237 411 252 417
rect 228 405 252 411
rect 228 399 231 405
rect 237 399 252 405
rect 228 396 252 399
rect -324 381 -312 384
rect -324 375 -321 381
rect -315 375 -312 381
rect -348 333 -336 336
rect -348 327 -345 333
rect -339 327 -336 333
rect -348 285 -336 327
rect -348 279 -345 285
rect -339 279 -336 285
rect -348 237 -336 279
rect -348 231 -345 237
rect -339 231 -336 237
rect -348 189 -336 231
rect -348 183 -345 189
rect -339 183 -336 189
rect -348 45 -336 183
rect -348 39 -345 45
rect -339 39 -336 45
rect -348 33 -336 39
rect -348 27 -345 33
rect -339 27 -336 33
rect -348 21 -336 27
rect -348 15 -345 21
rect -339 15 -336 21
rect -348 -3 -336 15
rect -324 45 -312 375
rect -276 381 -264 396
rect -276 375 -273 381
rect -267 375 -264 381
rect -276 357 -264 375
rect -228 381 -216 384
rect -228 375 -225 381
rect -219 375 -216 381
rect -228 372 -216 375
rect -276 351 -273 357
rect -267 351 -264 357
rect -300 333 -288 336
rect -300 327 -297 333
rect -291 327 -288 333
rect -300 324 -288 327
rect -276 69 -264 351
rect -276 63 -273 69
rect -267 63 -264 69
rect -276 60 -264 63
rect -228 93 -216 96
rect -228 87 -225 93
rect -219 87 -216 93
rect -228 69 -216 87
rect -228 63 -225 69
rect -219 63 -216 69
rect -228 48 -216 63
rect -324 39 -321 45
rect -315 39 -312 45
rect -324 33 -312 39
rect -324 27 -321 33
rect -315 27 -312 33
rect -324 21 -312 27
rect -324 15 -321 21
rect -315 15 -312 21
rect -324 12 -312 15
rect -300 45 -288 48
rect -300 39 -297 45
rect -291 39 -288 45
rect -300 33 -288 39
rect -300 27 -297 33
rect -291 27 -288 33
rect -300 21 -288 27
rect -300 15 -297 21
rect -291 15 -288 21
rect -348 -9 -345 -3
rect -339 -9 -336 -3
rect -348 -12 -336 -9
rect -300 -3 -288 15
rect -276 45 -216 48
rect -276 39 -273 45
rect -267 39 -216 45
rect -276 36 -216 39
rect -204 45 -192 396
rect -180 381 -168 384
rect -180 375 -177 381
rect -171 375 -168 381
rect -180 372 -168 375
rect -132 381 -120 384
rect -132 375 -129 381
rect -123 375 -120 381
rect -132 357 -120 375
rect -84 381 -72 384
rect -84 375 -81 381
rect -75 375 -72 381
rect -84 372 -72 375
rect -132 351 -129 357
rect -123 351 -120 357
rect -132 348 -120 351
rect -156 333 -144 336
rect -156 327 -153 333
rect -147 327 -144 333
rect -156 309 -144 327
rect -156 303 -153 309
rect -147 303 -144 309
rect -156 285 -144 303
rect -156 279 -153 285
rect -147 279 -144 285
rect -156 237 -144 279
rect -156 231 -153 237
rect -147 231 -144 237
rect -156 189 -144 231
rect -156 183 -153 189
rect -147 183 -144 189
rect -156 141 -144 183
rect -156 135 -153 141
rect -147 135 -144 141
rect -180 93 -168 96
rect -180 87 -177 93
rect -171 87 -168 93
rect -180 69 -168 87
rect -180 63 -177 69
rect -171 63 -168 69
rect -180 60 -168 63
rect -204 39 -201 45
rect -195 39 -192 45
rect -276 33 -264 36
rect -276 27 -273 33
rect -267 27 -264 33
rect -276 21 -264 27
rect -204 33 -192 39
rect -204 27 -201 33
rect -195 27 -192 33
rect -276 15 -273 21
rect -267 15 -264 21
rect -276 12 -264 15
rect -252 21 -240 24
rect -252 15 -249 21
rect -243 15 -240 21
rect -300 -9 -297 -3
rect -291 -9 -288 -3
rect -300 -12 -288 -9
rect -252 -3 -240 15
rect -204 21 -192 27
rect -204 15 -201 21
rect -195 15 -192 21
rect -204 12 -192 15
rect -156 45 -144 135
rect -108 333 -96 336
rect -108 327 -105 333
rect -99 327 -96 333
rect -108 285 -96 327
rect -108 279 -105 285
rect -99 279 -96 285
rect -108 237 -96 279
rect -108 231 -105 237
rect -99 231 -96 237
rect -108 189 -96 231
rect -108 183 -105 189
rect -99 183 -96 189
rect -108 141 -96 183
rect -108 135 -105 141
rect -99 135 -96 141
rect -132 93 -120 96
rect -132 87 -129 93
rect -123 87 -120 93
rect -132 69 -120 87
rect -132 63 -129 69
rect -123 63 -120 69
rect -132 60 -120 63
rect -156 39 -153 45
rect -147 39 -144 45
rect -156 33 -144 39
rect -156 27 -153 33
rect -147 27 -144 33
rect -156 21 -144 27
rect -156 15 -153 21
rect -147 15 -144 21
rect -252 -9 -249 -3
rect -243 -9 -240 -3
rect -252 -12 -240 -9
rect -156 -3 -144 15
rect -156 -9 -153 -3
rect -147 -9 -144 -3
rect -156 -12 -144 -9
rect -108 45 -96 135
rect -60 261 -48 396
rect -36 381 -24 384
rect -36 375 -33 381
rect -27 375 -24 381
rect -36 372 -24 375
rect 12 381 24 384
rect 12 375 15 381
rect 21 375 24 381
rect 12 372 24 375
rect -60 255 -57 261
rect -51 255 -48 261
rect -84 69 -72 72
rect -84 63 -81 69
rect -75 63 -72 69
rect -84 60 -72 63
rect -108 39 -105 45
rect -99 39 -96 45
rect -108 33 -96 39
rect -108 27 -105 33
rect -99 27 -96 33
rect -108 21 -96 27
rect -108 15 -105 21
rect -99 15 -96 21
rect -108 -3 -96 15
rect -60 45 -48 255
rect -12 333 0 336
rect -12 327 -9 333
rect -3 327 0 333
rect -12 285 0 327
rect -12 279 -9 285
rect -3 279 0 285
rect -12 237 0 279
rect -12 231 -9 237
rect -3 231 0 237
rect -12 189 0 231
rect -12 183 -9 189
rect -3 183 0 189
rect -36 69 -24 72
rect -36 63 -33 69
rect -27 63 -24 69
rect -36 60 -24 63
rect -60 39 -57 45
rect -51 39 -48 45
rect -60 33 -48 39
rect -60 27 -57 33
rect -51 27 -48 33
rect -60 21 -48 27
rect -60 15 -57 21
rect -51 15 -48 21
rect -60 12 -48 15
rect -12 45 0 183
rect 36 117 48 396
rect 60 381 72 384
rect 60 375 63 381
rect 69 375 72 381
rect 60 372 72 375
rect 108 381 120 384
rect 108 375 111 381
rect 117 375 120 381
rect 108 357 120 375
rect 108 351 111 357
rect 117 351 120 357
rect 108 348 120 351
rect 156 381 168 384
rect 156 375 159 381
rect 165 375 168 381
rect 156 357 168 375
rect 156 351 159 357
rect 165 351 168 357
rect 156 348 168 351
rect 204 381 216 384
rect 204 375 207 381
rect 213 375 216 381
rect 204 357 216 375
rect 204 351 207 357
rect 213 351 216 357
rect 204 348 216 351
rect 36 111 39 117
rect 45 111 48 117
rect 12 69 24 72
rect 12 63 15 69
rect 21 63 24 69
rect 12 60 24 63
rect -12 39 -9 45
rect -3 39 0 45
rect -12 33 0 39
rect -12 27 -9 33
rect -3 27 0 33
rect -12 21 0 27
rect -12 15 -9 21
rect -3 15 0 21
rect -108 -9 -105 -3
rect -99 -9 -96 -3
rect -108 -12 -96 -9
rect -12 -3 0 15
rect 36 45 48 111
rect 84 333 96 336
rect 84 327 87 333
rect 93 327 96 333
rect 84 285 96 327
rect 84 279 87 285
rect 93 279 96 285
rect 84 237 96 279
rect 84 231 87 237
rect 93 231 96 237
rect 84 189 96 231
rect 84 183 87 189
rect 93 183 96 189
rect 60 69 72 72
rect 60 63 63 69
rect 69 63 72 69
rect 60 60 72 63
rect 36 39 39 45
rect 45 39 48 45
rect 36 33 48 39
rect 36 27 39 33
rect 45 27 48 33
rect 36 21 48 27
rect 36 15 39 21
rect 45 15 48 21
rect 36 12 48 15
rect 84 45 96 183
rect 180 333 192 336
rect 180 327 183 333
rect 189 327 192 333
rect 180 285 192 327
rect 180 279 183 285
rect 189 279 192 285
rect 180 237 192 279
rect 180 231 183 237
rect 189 231 192 237
rect 180 189 192 231
rect 180 183 183 189
rect 189 183 192 189
rect 132 165 144 168
rect 132 159 135 165
rect 141 159 144 165
rect 108 69 120 72
rect 108 63 111 69
rect 117 63 120 69
rect 108 60 120 63
rect 84 39 87 45
rect 93 39 96 45
rect 84 33 96 39
rect 84 27 87 33
rect 93 27 96 33
rect 84 21 96 27
rect 84 15 87 21
rect 93 15 96 21
rect -12 -9 -9 -3
rect -3 -9 0 -3
rect -12 -12 0 -9
rect 84 -3 96 15
rect 132 45 144 159
rect 156 69 168 72
rect 156 63 159 69
rect 165 63 168 69
rect 156 60 168 63
rect 132 39 135 45
rect 141 39 144 45
rect 132 33 144 39
rect 132 27 135 33
rect 141 27 144 33
rect 132 21 144 27
rect 132 15 135 21
rect 141 15 144 21
rect 132 12 144 15
rect 180 45 192 183
rect 228 333 240 336
rect 228 327 231 333
rect 237 327 240 333
rect 228 285 240 327
rect 228 279 231 285
rect 237 279 240 285
rect 228 237 240 279
rect 228 231 231 237
rect 237 231 240 237
rect 228 189 240 231
rect 228 183 231 189
rect 237 183 240 189
rect 204 93 216 96
rect 204 87 207 93
rect 213 87 216 93
rect 204 69 216 87
rect 204 63 207 69
rect 213 63 216 69
rect 204 60 216 63
rect 180 39 183 45
rect 189 39 192 45
rect 180 33 192 39
rect 180 27 183 33
rect 189 27 192 33
rect 180 21 192 27
rect 180 15 183 21
rect 189 15 192 21
rect 84 -9 87 -3
rect 93 -9 96 -3
rect 84 -12 96 -9
rect 180 -3 192 15
rect 180 -9 183 -3
rect 189 -9 192 -3
rect 180 -12 192 -9
rect 228 45 240 183
rect 228 39 231 45
rect 237 39 240 45
rect 228 33 240 39
rect 228 27 231 33
rect 237 27 240 33
rect 228 21 240 27
rect 228 15 231 21
rect 237 15 240 21
rect 228 -3 240 15
rect 228 -9 231 -3
rect 237 -9 240 -3
rect 228 -12 240 -9
<< via2 >>
rect -321 567 -315 573
rect -273 567 -267 573
rect -225 567 -219 573
rect -177 567 -171 573
rect -129 567 -123 573
rect -81 567 -75 573
rect -33 567 -27 573
rect 15 567 21 573
rect 63 567 69 573
rect 111 567 117 573
rect 159 567 165 573
rect 207 567 213 573
rect -345 543 -339 549
rect -345 531 -339 537
rect -345 519 -339 525
rect -345 495 -339 501
rect -297 543 -291 549
rect -297 531 -291 537
rect -297 519 -291 525
rect -321 471 -315 477
rect -249 543 -243 549
rect -249 531 -243 537
rect -249 519 -243 525
rect -273 471 -267 477
rect -201 543 -195 549
rect -201 531 -195 537
rect -201 519 -195 525
rect -225 447 -219 453
rect -153 543 -147 549
rect -153 531 -147 537
rect -153 519 -147 525
rect -177 447 -171 453
rect -105 543 -99 549
rect -105 531 -99 537
rect -105 519 -99 525
rect -129 471 -123 477
rect -57 543 -51 549
rect -57 531 -51 537
rect -57 519 -51 525
rect -81 471 -75 477
rect -9 543 -3 549
rect -9 531 -3 537
rect -9 519 -3 525
rect -33 471 -27 477
rect 39 543 45 549
rect 39 531 45 537
rect 39 519 45 525
rect 15 471 21 477
rect 87 543 93 549
rect 87 531 93 537
rect 87 519 93 525
rect 63 471 69 477
rect 135 543 141 549
rect 135 531 141 537
rect 135 519 141 525
rect 111 471 117 477
rect 183 543 189 549
rect 183 531 189 537
rect 183 519 189 525
rect 159 471 165 477
rect 231 543 237 549
rect 231 531 237 537
rect 231 519 237 525
rect 207 471 213 477
rect -105 423 -99 429
rect -57 423 -51 429
rect -9 423 -3 429
rect 39 423 45 429
rect 87 423 93 429
rect 135 423 141 429
rect 183 423 189 429
rect 231 423 237 429
rect -105 411 -99 417
rect -9 411 -3 417
rect -105 399 -99 405
rect 87 411 93 417
rect -9 399 -3 405
rect 87 399 93 405
rect 135 411 141 417
rect 135 399 141 405
rect 183 411 189 417
rect 183 399 189 405
rect 231 411 237 417
rect 231 399 237 405
rect -345 327 -339 333
rect -345 279 -339 285
rect -345 231 -339 237
rect -345 183 -339 189
rect -345 39 -339 45
rect -345 27 -339 33
rect -345 15 -339 21
rect -225 375 -219 381
rect -273 351 -267 357
rect -297 327 -291 333
rect -225 87 -219 93
rect -297 39 -291 45
rect -297 27 -291 33
rect -297 15 -291 21
rect -177 375 -171 381
rect -81 375 -75 381
rect -129 351 -123 357
rect -153 327 -147 333
rect -153 303 -147 309
rect -153 279 -147 285
rect -153 231 -147 237
rect -153 183 -147 189
rect -153 135 -147 141
rect -177 87 -171 93
rect -201 39 -195 45
rect -201 27 -195 33
rect -249 15 -243 21
rect -201 15 -195 21
rect -105 327 -99 333
rect -105 279 -99 285
rect -105 231 -99 237
rect -105 183 -99 189
rect -105 135 -99 141
rect -129 87 -123 93
rect -153 39 -147 45
rect -153 27 -147 33
rect -153 15 -147 21
rect -33 375 -27 381
rect 15 375 21 381
rect -57 255 -51 261
rect -81 63 -75 69
rect -105 39 -99 45
rect -105 27 -99 33
rect -105 15 -99 21
rect -9 327 -3 333
rect -9 279 -3 285
rect -9 231 -3 237
rect -9 183 -3 189
rect -33 63 -27 69
rect 63 375 69 381
rect 111 351 117 357
rect 159 351 165 357
rect 207 351 213 357
rect 39 111 45 117
rect 15 63 21 69
rect -9 39 -3 45
rect -9 27 -3 33
rect -9 15 -3 21
rect 87 327 93 333
rect 87 279 93 285
rect 87 231 93 237
rect 87 183 93 189
rect 63 63 69 69
rect 183 327 189 333
rect 183 279 189 285
rect 183 231 189 237
rect 183 183 189 189
rect 135 159 141 165
rect 111 63 117 69
rect 87 39 93 45
rect 87 27 93 33
rect 87 15 93 21
rect 159 63 165 69
rect 231 327 237 333
rect 231 279 237 285
rect 231 231 237 237
rect 231 183 237 189
rect 207 87 213 93
rect 183 39 189 45
rect 183 27 189 33
rect 183 15 189 21
rect 231 39 237 45
rect 231 27 237 33
rect 231 15 237 21
<< metal3 >>
rect -396 573 288 576
rect -396 567 -321 573
rect -315 567 -273 573
rect -267 567 -225 573
rect -219 567 -177 573
rect -171 567 -129 573
rect -123 567 -81 573
rect -75 567 -33 573
rect -27 567 15 573
rect 21 567 63 573
rect 69 567 111 573
rect 117 567 159 573
rect 165 567 207 573
rect 213 567 288 573
rect -396 564 288 567
rect -396 549 288 552
rect -396 543 -345 549
rect -339 543 -297 549
rect -291 543 -249 549
rect -243 543 -201 549
rect -195 543 -153 549
rect -147 543 -105 549
rect -99 543 -57 549
rect -51 543 -9 549
rect -3 543 39 549
rect 45 543 87 549
rect 93 543 135 549
rect 141 543 183 549
rect 189 543 231 549
rect 237 543 288 549
rect -396 537 288 543
rect -396 531 -345 537
rect -339 531 -297 537
rect -291 531 -249 537
rect -243 531 -201 537
rect -195 531 -153 537
rect -147 531 -105 537
rect -99 531 -57 537
rect -51 531 -9 537
rect -3 531 39 537
rect 45 531 87 537
rect 93 531 135 537
rect 141 531 183 537
rect 189 531 231 537
rect 237 531 288 537
rect -396 525 288 531
rect -396 519 -345 525
rect -339 519 -297 525
rect -291 519 -249 525
rect -243 519 -201 525
rect -195 519 -153 525
rect -147 519 -105 525
rect -99 519 -57 525
rect -51 519 -9 525
rect -3 519 39 525
rect 45 519 87 525
rect 93 519 135 525
rect 141 519 183 525
rect 189 519 231 525
rect 237 519 288 525
rect -396 516 288 519
rect -372 504 -360 516
rect 252 504 264 516
rect -372 501 264 504
rect -372 495 -345 501
rect -339 495 264 501
rect -372 492 264 495
rect -396 477 288 480
rect -396 471 -321 477
rect -315 471 -273 477
rect -267 471 -129 477
rect -123 471 -81 477
rect -75 471 -33 477
rect -27 471 15 477
rect 21 471 63 477
rect 69 471 111 477
rect 117 471 159 477
rect 165 471 207 477
rect 213 471 288 477
rect -396 468 288 471
rect -396 453 288 456
rect -396 447 -225 453
rect -219 447 -177 453
rect -171 447 288 453
rect -396 444 288 447
rect -396 429 288 432
rect -396 423 -105 429
rect -99 423 -57 429
rect -51 423 -9 429
rect -3 423 39 429
rect 45 423 87 429
rect 93 423 135 429
rect 141 423 183 429
rect 189 423 231 429
rect 237 423 288 429
rect -396 417 288 423
rect -396 411 -105 417
rect -99 411 -9 417
rect -3 411 87 417
rect 93 411 135 417
rect 141 411 183 417
rect 189 411 231 417
rect 237 411 288 417
rect -396 405 288 411
rect -396 399 -105 405
rect -99 399 -9 405
rect -3 399 87 405
rect 93 399 135 405
rect 141 399 183 405
rect 189 399 231 405
rect 237 399 288 405
rect -396 396 288 399
rect -228 381 -216 384
rect -228 375 -225 381
rect -219 375 -216 381
rect -228 372 -216 375
rect -180 381 -168 384
rect -180 375 -177 381
rect -171 375 -168 381
rect -180 372 -168 375
rect -84 381 -72 384
rect -84 375 -81 381
rect -75 375 -72 381
rect -84 372 -72 375
rect -36 381 -24 384
rect -36 375 -33 381
rect -27 375 -24 381
rect -36 372 -24 375
rect 12 381 24 384
rect 12 375 15 381
rect 21 375 24 381
rect 12 372 24 375
rect 60 381 72 384
rect 60 375 63 381
rect 69 375 72 381
rect 60 372 72 375
rect -372 357 264 360
rect -372 351 -273 357
rect -267 351 -129 357
rect -123 351 111 357
rect 117 351 159 357
rect 165 351 207 357
rect 213 351 264 357
rect -372 348 264 351
rect -396 333 288 336
rect -396 327 -345 333
rect -339 327 -297 333
rect -291 327 -153 333
rect -147 327 -105 333
rect -99 327 -9 333
rect -3 327 87 333
rect 93 327 183 333
rect 189 327 231 333
rect 237 327 288 333
rect -396 324 288 327
rect -348 309 240 312
rect -348 303 -153 309
rect -147 303 240 309
rect -348 300 240 303
rect -348 285 240 288
rect -348 279 -345 285
rect -339 279 -153 285
rect -147 279 -105 285
rect -99 279 -9 285
rect -3 279 87 285
rect 93 279 183 285
rect 189 279 231 285
rect 237 279 240 285
rect -348 276 240 279
rect -348 261 252 264
rect -348 255 -225 261
rect -219 255 -177 261
rect -171 255 -57 261
rect -51 255 252 261
rect -348 252 252 255
rect -348 237 240 240
rect -348 231 -345 237
rect -339 231 -153 237
rect -147 231 -105 237
rect -99 231 -9 237
rect -3 231 87 237
rect 93 231 183 237
rect 189 231 231 237
rect 237 231 240 237
rect -348 228 240 231
rect -360 213 240 216
rect -360 207 -81 213
rect -75 207 -33 213
rect -27 207 240 213
rect -360 204 240 207
rect -348 189 240 192
rect -348 183 -345 189
rect -339 183 -153 189
rect -147 183 -105 189
rect -99 183 -9 189
rect -3 183 87 189
rect 93 183 183 189
rect 189 183 231 189
rect 237 183 240 189
rect -348 180 240 183
rect -348 165 252 168
rect -348 159 135 165
rect 141 159 252 165
rect -348 156 252 159
rect -348 141 240 144
rect -348 135 -153 141
rect -147 135 -105 141
rect -99 135 240 141
rect -348 132 240 135
rect -348 117 252 120
rect -348 111 15 117
rect 21 111 39 117
rect 45 111 63 117
rect 69 111 111 117
rect 117 111 159 117
rect 165 111 252 117
rect -348 108 252 111
rect -348 93 240 96
rect -348 87 -225 93
rect -219 87 -177 93
rect -171 87 -129 93
rect -123 87 207 93
rect 213 87 240 93
rect -348 84 240 87
rect -84 69 -72 72
rect -84 63 -81 69
rect -75 63 -72 69
rect -84 60 -72 63
rect -36 69 -24 72
rect -36 63 -33 69
rect -27 63 -24 69
rect -36 60 -24 63
rect 12 69 24 72
rect 12 63 15 69
rect 21 63 24 69
rect 12 60 24 63
rect 60 69 72 72
rect 60 63 63 69
rect 69 63 72 69
rect 60 60 72 63
rect 108 69 120 72
rect 108 63 111 69
rect 117 63 120 69
rect 108 60 120 63
rect 156 69 168 72
rect 156 63 159 69
rect 165 63 168 69
rect 156 60 168 63
rect -396 45 288 48
rect -396 39 -345 45
rect -339 39 -297 45
rect -291 39 -201 45
rect -195 39 -153 45
rect -147 39 -105 45
rect -99 39 -9 45
rect -3 39 87 45
rect 93 39 183 45
rect 189 39 231 45
rect 237 39 288 45
rect -396 33 288 39
rect -396 27 -345 33
rect -339 27 -297 33
rect -291 27 -201 33
rect -195 27 -153 33
rect -147 27 -105 33
rect -99 27 -9 33
rect -3 27 87 33
rect 93 27 183 33
rect 189 27 231 33
rect 237 27 288 33
rect -396 21 288 27
rect -396 15 -345 21
rect -339 15 -297 21
rect -291 15 -249 21
rect -243 15 -201 21
rect -195 15 -153 21
rect -147 15 -105 21
rect -99 15 -9 21
rect -3 15 87 21
rect 93 15 183 21
rect 189 15 231 21
rect 237 15 288 21
rect -396 12 288 15
<< via3 >>
rect -225 375 -219 381
rect -177 375 -171 381
rect -81 375 -75 381
rect -33 375 -27 381
rect 15 375 21 381
rect 63 375 69 381
rect -225 255 -219 261
rect -177 255 -171 261
rect -81 207 -75 213
rect -33 207 -27 213
rect 15 111 21 117
rect 63 111 69 117
rect 111 111 117 117
rect 159 111 165 117
rect -81 63 -75 69
rect -33 63 -27 69
rect 15 63 21 69
rect 63 63 69 69
rect 111 63 117 69
rect 159 63 165 69
<< metal4 >>
rect -228 381 -216 384
rect -228 375 -225 381
rect -219 375 -216 381
rect -228 372 -216 375
rect -180 381 -168 384
rect -180 375 -177 381
rect -171 375 -168 381
rect -180 372 -168 375
rect -84 381 -72 384
rect -84 375 -81 381
rect -75 375 -72 381
rect -84 372 -72 375
rect -36 381 -24 384
rect -36 375 -33 381
rect -27 375 -24 381
rect -36 372 -24 375
rect 12 381 24 384
rect 12 375 15 381
rect 21 375 24 381
rect 12 372 24 375
rect 60 381 72 384
rect 60 375 63 381
rect 69 375 72 381
rect 60 372 72 375
rect -228 261 -216 264
rect -228 255 -225 261
rect -219 255 -216 261
rect -228 252 -216 255
rect -180 261 -168 264
rect -180 255 -177 261
rect -171 255 -168 261
rect -180 252 -168 255
rect -84 213 -72 216
rect -84 207 -81 213
rect -75 207 -72 213
rect -84 204 -72 207
rect -36 213 -24 216
rect -36 207 -33 213
rect -27 207 -24 213
rect -36 204 -24 207
rect 12 117 24 120
rect 12 111 15 117
rect 21 111 24 117
rect 12 108 24 111
rect 60 117 72 120
rect 60 111 63 117
rect 69 111 72 117
rect 60 108 72 111
rect 108 117 120 120
rect 108 111 111 117
rect 117 111 120 117
rect 108 108 120 111
rect 156 117 168 120
rect 156 111 159 117
rect 165 111 168 117
rect 156 108 168 111
rect -84 69 -72 72
rect -84 63 -81 69
rect -75 63 -72 69
rect -84 60 -72 63
rect -36 69 -24 72
rect -36 63 -33 69
rect -27 63 -24 69
rect -36 60 -24 63
rect 12 69 24 72
rect 12 63 15 69
rect 21 63 24 69
rect 12 60 24 63
rect 60 69 72 72
rect 60 63 63 69
rect 69 63 72 69
rect 60 60 72 63
rect 108 69 120 72
rect 108 63 111 69
rect 117 63 120 69
rect 108 60 120 63
rect 156 69 168 72
rect 156 63 159 69
rect 165 63 168 69
rect 156 60 168 63
<< via4 >>
rect -225 375 -219 381
rect -177 375 -171 381
rect -81 375 -75 381
rect -33 375 -27 381
rect 15 375 21 381
rect 63 375 69 381
rect -225 255 -219 261
rect -177 255 -171 261
rect -81 207 -75 213
rect -33 207 -27 213
rect 15 111 21 117
rect 63 111 69 117
rect 111 111 117 117
rect 159 111 165 117
rect -81 63 -75 69
rect -33 63 -27 69
rect 15 63 21 69
rect 63 63 69 69
rect 111 63 117 69
rect 159 63 165 69
<< metal5 >>
rect -228 381 -216 384
rect -228 375 -225 381
rect -219 375 -216 381
rect -228 261 -216 375
rect -228 255 -225 261
rect -219 255 -216 261
rect -228 252 -216 255
rect -180 381 -168 384
rect -180 375 -177 381
rect -171 375 -168 381
rect -180 261 -168 375
rect -180 255 -177 261
rect -171 255 -168 261
rect -180 252 -168 255
rect -84 381 -72 384
rect -84 375 -81 381
rect -75 375 -72 381
rect -84 213 -72 375
rect -84 207 -81 213
rect -75 207 -72 213
rect -84 69 -72 207
rect -84 63 -81 69
rect -75 63 -72 69
rect -84 60 -72 63
rect -36 381 -24 384
rect -36 375 -33 381
rect -27 375 -24 381
rect -36 213 -24 375
rect -36 207 -33 213
rect -27 207 -24 213
rect -36 69 -24 207
rect -36 63 -33 69
rect -27 63 -24 69
rect -36 60 -24 63
rect 12 381 24 384
rect 12 375 15 381
rect 21 375 24 381
rect 12 117 24 375
rect 12 111 15 117
rect 21 111 24 117
rect 12 69 24 111
rect 12 63 15 69
rect 21 63 24 69
rect 12 60 24 63
rect 60 381 72 384
rect 60 375 63 381
rect 69 375 72 381
rect 60 117 72 375
rect 60 111 63 117
rect 69 111 72 117
rect 60 69 72 111
rect 60 63 63 69
rect 69 63 72 69
rect 60 60 72 63
rect 108 117 120 120
rect 108 111 111 117
rect 117 111 120 117
rect 108 69 120 111
rect 108 63 111 69
rect 117 63 120 69
rect 108 60 120 63
rect 156 117 168 120
rect 156 111 159 117
rect 165 111 168 117
rect 156 69 168 111
rect 156 63 159 69
rect 165 63 168 69
rect 156 60 168 63
<< labels >>
rlabel metal3 -360 204 -348 216 0 ref
port 1 nsew
rlabel metal3 240 156 252 168 0 iq
port 2 nsew
rlabel metal3 -396 516 288 552 0 vhi
port 3 nsew
rlabel metal3 -396 396 288 432 0 vdd
port 5 nsew
rlabel metal3 -396 444 288 456 0 bp
port 6 nsew
rlabel metal3 -396 12 288 48 0 vss
port 7 nsew
rlabel metal3 240 108 252 120 0 q
rlabel metal3 240 252 252 264 0 x
rlabel metal2 -228 72 -216 84 0 vlo
rlabel metal3 -396 564 288 576 0 gp
port 4 nsew
rlabel metal3 -276 348 -264 360 0 tihi
<< end >>
