magic
tech gf180mcuC
timestamp 1697225838
<< nwell >>
rect -42 342 1518 606
<< nmos >>
rect 0 12 12 48
rect 24 12 36 48
rect 48 12 60 48
rect 72 12 84 48
rect 96 12 108 48
rect 120 12 132 48
rect 144 12 156 48
rect 168 12 180 48
rect 216 12 228 48
rect 240 12 252 48
rect 264 12 276 48
rect 288 12 300 48
rect 312 12 324 48
rect 336 12 348 48
rect 360 12 372 48
rect 384 12 396 48
rect 432 12 444 48
rect 456 12 468 48
rect 480 12 492 48
rect 504 12 516 48
rect 528 12 540 48
rect 552 12 564 48
rect 576 12 588 48
rect 600 12 612 48
rect 648 12 660 48
rect 672 12 684 48
rect 696 12 708 48
rect 720 12 732 48
rect 744 12 756 48
rect 768 12 780 48
rect 792 12 804 48
rect 816 12 828 48
rect 864 12 876 48
rect 888 12 900 48
rect 912 12 924 48
rect 936 12 948 48
rect 960 12 972 48
rect 984 12 996 48
rect 1008 12 1020 48
rect 1032 12 1044 48
rect 1080 12 1092 48
rect 1104 12 1116 48
rect 1128 12 1140 48
rect 1152 12 1164 48
rect 1176 12 1188 48
rect 1200 12 1212 48
rect 1224 12 1236 48
rect 1248 12 1260 48
rect 1296 12 1308 48
rect 1320 12 1332 48
rect 1344 12 1356 48
rect 1368 12 1380 48
rect 1392 12 1404 48
rect 1416 12 1428 48
rect 1440 12 1452 48
rect 1464 12 1476 48
<< mvnmos >>
rect 0 252 12 288
rect 24 252 36 288
rect 48 252 60 288
rect 72 252 84 288
rect 96 252 108 288
rect 120 252 132 288
rect 144 252 156 288
rect 168 252 180 288
rect 216 252 228 288
rect 240 252 252 288
rect 264 252 276 288
rect 288 252 300 288
rect 312 252 324 288
rect 336 252 348 288
rect 360 252 372 288
rect 384 252 396 288
rect 432 252 444 288
rect 456 252 468 288
rect 480 252 492 288
rect 504 252 516 288
rect 528 252 540 288
rect 552 252 564 288
rect 576 252 588 288
rect 600 252 612 288
rect 648 252 660 288
rect 672 252 684 288
rect 696 252 708 288
rect 720 252 732 288
rect 744 252 756 288
rect 768 252 780 288
rect 792 252 804 288
rect 816 252 828 288
rect 864 252 876 288
rect 912 252 924 288
rect 936 252 948 288
rect 960 252 972 288
rect 984 252 996 288
rect 1008 252 1020 288
rect 1032 252 1044 288
rect 1080 252 1092 288
rect 1104 252 1116 288
rect 1128 252 1140 288
rect 1152 252 1164 288
rect 1176 252 1188 288
rect 1200 252 1212 288
rect 1224 252 1236 288
rect 1248 252 1260 288
rect 1296 252 1308 288
rect 1320 252 1332 288
rect 1344 252 1356 288
rect 1368 252 1380 288
rect 1392 252 1404 288
rect 1416 252 1428 288
rect 1440 252 1452 288
rect 1464 252 1476 288
<< mvpmos >>
rect 0 540 12 576
rect 24 540 36 576
rect 48 540 60 576
rect 72 540 84 576
rect 96 540 108 576
rect 120 540 132 576
rect 144 540 156 576
rect 168 540 180 576
rect 216 540 228 576
rect 240 540 252 576
rect 264 540 276 576
rect 288 540 300 576
rect 312 540 324 576
rect 336 540 348 576
rect 360 540 372 576
rect 384 540 396 576
rect 432 540 444 576
rect 456 540 468 576
rect 480 540 492 576
rect 504 540 516 576
rect 528 540 540 576
rect 552 540 564 576
rect 576 540 588 576
rect 600 540 612 576
rect 648 540 660 576
rect 672 540 684 576
rect 696 540 708 576
rect 720 540 732 576
rect 744 540 756 576
rect 768 540 780 576
rect 792 540 804 576
rect 816 540 828 576
rect 864 540 876 576
rect 888 540 900 576
rect 912 540 924 576
rect 936 540 948 576
rect 960 540 972 576
rect 984 540 996 576
rect 1008 540 1020 576
rect 1032 540 1044 576
rect 1080 540 1092 576
rect 1104 540 1116 576
rect 1128 540 1140 576
rect 1152 540 1164 576
rect 1176 540 1188 576
rect 1200 540 1212 576
rect 1224 540 1236 576
rect 1248 540 1260 576
rect 1296 540 1308 576
rect 1320 540 1332 576
rect 1344 540 1356 576
rect 1368 540 1380 576
rect 1392 540 1404 576
rect 1416 540 1428 576
rect 1440 540 1452 576
rect 1464 540 1476 576
rect 0 444 12 480
rect 24 444 36 480
rect 48 444 60 480
rect 72 444 84 480
rect 96 444 108 480
rect 120 444 132 480
rect 144 444 156 480
rect 168 444 180 480
rect 216 444 228 480
rect 240 444 252 480
rect 264 444 276 480
rect 288 444 300 480
rect 312 444 324 480
rect 336 444 348 480
rect 360 444 372 480
rect 384 444 396 480
rect 432 444 444 480
rect 456 444 468 480
rect 480 444 492 480
rect 504 444 516 480
rect 528 444 540 480
rect 552 444 564 480
rect 576 444 588 480
rect 600 444 612 480
rect 648 444 660 480
rect 672 444 684 480
rect 696 444 708 480
rect 720 444 732 480
rect 744 444 756 480
rect 768 444 780 480
rect 792 444 804 480
rect 816 444 828 480
rect 864 444 876 480
rect 888 444 900 480
rect 912 444 924 480
rect 936 444 948 480
rect 960 444 972 480
rect 984 444 996 480
rect 1008 444 1020 480
rect 1032 444 1044 480
rect 1080 444 1092 480
rect 1104 444 1116 480
rect 1128 444 1140 480
rect 1152 444 1164 480
rect 1176 444 1188 480
rect 1200 444 1212 480
rect 1224 444 1236 480
rect 1248 444 1260 480
rect 1296 444 1308 480
rect 1320 444 1332 480
rect 1344 444 1356 480
rect 1368 444 1380 480
rect 1392 444 1404 480
rect 1416 444 1428 480
rect 1440 444 1452 480
rect 1464 444 1476 480
<< ndiff >>
rect -12 45 0 48
rect -12 39 -9 45
rect -3 39 0 45
rect -12 33 0 39
rect -12 27 -9 33
rect -3 27 0 33
rect -12 21 0 27
rect -12 15 -9 21
rect -3 15 0 21
rect -12 12 0 15
rect 12 12 24 48
rect 36 45 48 48
rect 36 39 39 45
rect 45 39 48 45
rect 36 33 48 39
rect 36 27 39 33
rect 45 27 48 33
rect 36 21 48 27
rect 36 15 39 21
rect 45 15 48 21
rect 36 12 48 15
rect 60 12 72 48
rect 84 45 96 48
rect 84 39 87 45
rect 93 39 96 45
rect 84 33 96 39
rect 84 27 87 33
rect 93 27 96 33
rect 84 21 96 27
rect 84 15 87 21
rect 93 15 96 21
rect 84 12 96 15
rect 108 12 120 48
rect 132 45 144 48
rect 132 39 135 45
rect 141 39 144 45
rect 132 33 144 39
rect 132 27 135 33
rect 141 27 144 33
rect 132 21 144 27
rect 132 15 135 21
rect 141 15 144 21
rect 132 12 144 15
rect 156 12 168 48
rect 180 45 192 48
rect 180 39 183 45
rect 189 39 192 45
rect 180 33 192 39
rect 180 27 183 33
rect 189 27 192 33
rect 180 21 192 27
rect 180 15 183 21
rect 189 15 192 21
rect 180 12 192 15
rect 204 45 216 48
rect 204 39 207 45
rect 213 39 216 45
rect 204 33 216 39
rect 204 27 207 33
rect 213 27 216 33
rect 204 21 216 27
rect 204 15 207 21
rect 213 15 216 21
rect 204 12 216 15
rect 228 12 240 48
rect 252 45 264 48
rect 252 39 255 45
rect 261 39 264 45
rect 252 33 264 39
rect 252 27 255 33
rect 261 27 264 33
rect 252 21 264 27
rect 252 15 255 21
rect 261 15 264 21
rect 252 12 264 15
rect 276 12 288 48
rect 300 45 312 48
rect 300 39 303 45
rect 309 39 312 45
rect 300 33 312 39
rect 300 27 303 33
rect 309 27 312 33
rect 300 21 312 27
rect 300 15 303 21
rect 309 15 312 21
rect 300 12 312 15
rect 324 12 336 48
rect 348 45 360 48
rect 348 39 351 45
rect 357 39 360 45
rect 348 33 360 39
rect 348 27 351 33
rect 357 27 360 33
rect 348 21 360 27
rect 348 15 351 21
rect 357 15 360 21
rect 348 12 360 15
rect 372 12 384 48
rect 396 45 408 48
rect 396 39 399 45
rect 405 39 408 45
rect 396 33 408 39
rect 396 27 399 33
rect 405 27 408 33
rect 396 21 408 27
rect 396 15 399 21
rect 405 15 408 21
rect 396 12 408 15
rect 420 45 432 48
rect 420 39 423 45
rect 429 39 432 45
rect 420 33 432 39
rect 420 27 423 33
rect 429 27 432 33
rect 420 21 432 27
rect 420 15 423 21
rect 429 15 432 21
rect 420 12 432 15
rect 444 12 456 48
rect 468 12 480 48
rect 492 12 504 48
rect 516 45 528 48
rect 516 39 519 45
rect 525 39 528 45
rect 516 33 528 39
rect 516 27 519 33
rect 525 27 528 33
rect 516 21 528 27
rect 516 15 519 21
rect 525 15 528 21
rect 516 12 528 15
rect 540 12 552 48
rect 564 12 576 48
rect 588 12 600 48
rect 612 45 624 48
rect 612 39 615 45
rect 621 39 624 45
rect 612 33 624 39
rect 612 27 615 33
rect 621 27 624 33
rect 612 21 624 27
rect 612 15 615 21
rect 621 15 624 21
rect 612 12 624 15
rect 636 45 648 48
rect 636 39 639 45
rect 645 39 648 45
rect 636 33 648 39
rect 636 27 639 33
rect 645 27 648 33
rect 636 21 648 27
rect 636 15 639 21
rect 645 15 648 21
rect 636 12 648 15
rect 660 12 672 48
rect 684 12 696 48
rect 708 12 720 48
rect 732 45 744 48
rect 732 39 735 45
rect 741 39 744 45
rect 732 33 744 39
rect 732 27 735 33
rect 741 27 744 33
rect 732 21 744 27
rect 732 15 735 21
rect 741 15 744 21
rect 732 12 744 15
rect 756 12 768 48
rect 780 12 792 48
rect 804 12 816 48
rect 828 45 840 48
rect 828 39 831 45
rect 837 39 840 45
rect 828 33 840 39
rect 828 27 831 33
rect 837 27 840 33
rect 828 21 840 27
rect 828 15 831 21
rect 837 15 840 21
rect 828 12 840 15
rect 852 45 864 48
rect 852 39 855 45
rect 861 39 864 45
rect 852 33 864 39
rect 852 27 855 33
rect 861 27 864 33
rect 852 21 864 27
rect 852 15 855 21
rect 861 15 864 21
rect 852 12 864 15
rect 876 12 888 48
rect 900 12 912 48
rect 924 12 936 48
rect 948 12 960 48
rect 972 12 984 48
rect 996 12 1008 48
rect 1020 12 1032 48
rect 1044 45 1056 48
rect 1044 39 1047 45
rect 1053 39 1056 45
rect 1044 33 1056 39
rect 1044 27 1047 33
rect 1053 27 1056 33
rect 1044 21 1056 27
rect 1044 15 1047 21
rect 1053 15 1056 21
rect 1044 12 1056 15
rect 1068 45 1080 48
rect 1068 39 1071 45
rect 1077 39 1080 45
rect 1068 33 1080 39
rect 1068 27 1071 33
rect 1077 27 1080 33
rect 1068 21 1080 27
rect 1068 15 1071 21
rect 1077 15 1080 21
rect 1068 12 1080 15
rect 1092 45 1104 48
rect 1092 39 1095 45
rect 1101 39 1104 45
rect 1092 33 1104 39
rect 1092 27 1095 33
rect 1101 27 1104 33
rect 1092 21 1104 27
rect 1092 15 1095 21
rect 1101 15 1104 21
rect 1092 12 1104 15
rect 1116 45 1128 48
rect 1116 39 1119 45
rect 1125 39 1128 45
rect 1116 33 1128 39
rect 1116 27 1119 33
rect 1125 27 1128 33
rect 1116 21 1128 27
rect 1116 15 1119 21
rect 1125 15 1128 21
rect 1116 12 1128 15
rect 1140 45 1152 48
rect 1140 39 1143 45
rect 1149 39 1152 45
rect 1140 33 1152 39
rect 1140 27 1143 33
rect 1149 27 1152 33
rect 1140 21 1152 27
rect 1140 15 1143 21
rect 1149 15 1152 21
rect 1140 12 1152 15
rect 1164 45 1176 48
rect 1164 39 1167 45
rect 1173 39 1176 45
rect 1164 33 1176 39
rect 1164 27 1167 33
rect 1173 27 1176 33
rect 1164 21 1176 27
rect 1164 15 1167 21
rect 1173 15 1176 21
rect 1164 12 1176 15
rect 1188 45 1200 48
rect 1188 39 1191 45
rect 1197 39 1200 45
rect 1188 33 1200 39
rect 1188 27 1191 33
rect 1197 27 1200 33
rect 1188 21 1200 27
rect 1188 15 1191 21
rect 1197 15 1200 21
rect 1188 12 1200 15
rect 1212 45 1224 48
rect 1212 39 1215 45
rect 1221 39 1224 45
rect 1212 33 1224 39
rect 1212 27 1215 33
rect 1221 27 1224 33
rect 1212 21 1224 27
rect 1212 15 1215 21
rect 1221 15 1224 21
rect 1212 12 1224 15
rect 1236 45 1248 48
rect 1236 39 1239 45
rect 1245 39 1248 45
rect 1236 33 1248 39
rect 1236 27 1239 33
rect 1245 27 1248 33
rect 1236 21 1248 27
rect 1236 15 1239 21
rect 1245 15 1248 21
rect 1236 12 1248 15
rect 1260 45 1272 48
rect 1260 39 1263 45
rect 1269 39 1272 45
rect 1260 33 1272 39
rect 1260 27 1263 33
rect 1269 27 1272 33
rect 1260 21 1272 27
rect 1260 15 1263 21
rect 1269 15 1272 21
rect 1260 12 1272 15
rect 1284 45 1296 48
rect 1284 39 1287 45
rect 1293 39 1296 45
rect 1284 33 1296 39
rect 1284 27 1287 33
rect 1293 27 1296 33
rect 1284 21 1296 27
rect 1284 15 1287 21
rect 1293 15 1296 21
rect 1284 12 1296 15
rect 1308 45 1320 48
rect 1308 39 1311 45
rect 1317 39 1320 45
rect 1308 33 1320 39
rect 1308 27 1311 33
rect 1317 27 1320 33
rect 1308 21 1320 27
rect 1308 15 1311 21
rect 1317 15 1320 21
rect 1308 12 1320 15
rect 1332 45 1344 48
rect 1332 39 1335 45
rect 1341 39 1344 45
rect 1332 33 1344 39
rect 1332 27 1335 33
rect 1341 27 1344 33
rect 1332 21 1344 27
rect 1332 15 1335 21
rect 1341 15 1344 21
rect 1332 12 1344 15
rect 1356 45 1368 48
rect 1356 39 1359 45
rect 1365 39 1368 45
rect 1356 33 1368 39
rect 1356 27 1359 33
rect 1365 27 1368 33
rect 1356 21 1368 27
rect 1356 15 1359 21
rect 1365 15 1368 21
rect 1356 12 1368 15
rect 1380 45 1392 48
rect 1380 39 1383 45
rect 1389 39 1392 45
rect 1380 33 1392 39
rect 1380 27 1383 33
rect 1389 27 1392 33
rect 1380 21 1392 27
rect 1380 15 1383 21
rect 1389 15 1392 21
rect 1380 12 1392 15
rect 1404 45 1416 48
rect 1404 39 1407 45
rect 1413 39 1416 45
rect 1404 33 1416 39
rect 1404 27 1407 33
rect 1413 27 1416 33
rect 1404 21 1416 27
rect 1404 15 1407 21
rect 1413 15 1416 21
rect 1404 12 1416 15
rect 1428 45 1440 48
rect 1428 39 1431 45
rect 1437 39 1440 45
rect 1428 33 1440 39
rect 1428 27 1431 33
rect 1437 27 1440 33
rect 1428 21 1440 27
rect 1428 15 1431 21
rect 1437 15 1440 21
rect 1428 12 1440 15
rect 1452 45 1464 48
rect 1452 39 1455 45
rect 1461 39 1464 45
rect 1452 33 1464 39
rect 1452 27 1455 33
rect 1461 27 1464 33
rect 1452 21 1464 27
rect 1452 15 1455 21
rect 1461 15 1464 21
rect 1452 12 1464 15
rect 1476 45 1488 48
rect 1476 39 1479 45
rect 1485 39 1488 45
rect 1476 33 1488 39
rect 1476 27 1479 33
rect 1485 27 1488 33
rect 1476 21 1488 27
rect 1476 15 1479 21
rect 1485 15 1488 21
rect 1476 12 1488 15
<< mvndiff >>
rect -12 285 0 288
rect -12 279 -9 285
rect -3 279 0 285
rect -12 273 0 279
rect -12 267 -9 273
rect -3 267 0 273
rect -12 261 0 267
rect -12 255 -9 261
rect -3 255 0 261
rect -12 252 0 255
rect 12 285 24 288
rect 12 279 15 285
rect 21 279 24 285
rect 12 273 24 279
rect 12 267 15 273
rect 21 267 24 273
rect 12 261 24 267
rect 12 255 15 261
rect 21 255 24 261
rect 12 252 24 255
rect 36 285 48 288
rect 36 279 39 285
rect 45 279 48 285
rect 36 273 48 279
rect 36 267 39 273
rect 45 267 48 273
rect 36 261 48 267
rect 36 255 39 261
rect 45 255 48 261
rect 36 252 48 255
rect 60 285 72 288
rect 60 279 63 285
rect 69 279 72 285
rect 60 273 72 279
rect 60 267 63 273
rect 69 267 72 273
rect 60 261 72 267
rect 60 255 63 261
rect 69 255 72 261
rect 60 252 72 255
rect 84 285 96 288
rect 84 279 87 285
rect 93 279 96 285
rect 84 273 96 279
rect 84 267 87 273
rect 93 267 96 273
rect 84 261 96 267
rect 84 255 87 261
rect 93 255 96 261
rect 84 252 96 255
rect 108 285 120 288
rect 108 279 111 285
rect 117 279 120 285
rect 108 273 120 279
rect 108 267 111 273
rect 117 267 120 273
rect 108 261 120 267
rect 108 255 111 261
rect 117 255 120 261
rect 108 252 120 255
rect 132 285 144 288
rect 132 279 135 285
rect 141 279 144 285
rect 132 273 144 279
rect 132 267 135 273
rect 141 267 144 273
rect 132 261 144 267
rect 132 255 135 261
rect 141 255 144 261
rect 132 252 144 255
rect 156 285 168 288
rect 156 279 159 285
rect 165 279 168 285
rect 156 273 168 279
rect 156 267 159 273
rect 165 267 168 273
rect 156 261 168 267
rect 156 255 159 261
rect 165 255 168 261
rect 156 252 168 255
rect 180 285 192 288
rect 180 279 183 285
rect 189 279 192 285
rect 180 273 192 279
rect 180 267 183 273
rect 189 267 192 273
rect 180 261 192 267
rect 180 255 183 261
rect 189 255 192 261
rect 180 252 192 255
rect 204 285 216 288
rect 204 279 207 285
rect 213 279 216 285
rect 204 273 216 279
rect 204 267 207 273
rect 213 267 216 273
rect 204 261 216 267
rect 204 255 207 261
rect 213 255 216 261
rect 204 252 216 255
rect 228 252 240 288
rect 252 252 264 288
rect 276 252 288 288
rect 300 285 312 288
rect 300 279 303 285
rect 309 279 312 285
rect 300 273 312 279
rect 300 267 303 273
rect 309 267 312 273
rect 300 261 312 267
rect 300 255 303 261
rect 309 255 312 261
rect 300 252 312 255
rect 324 252 336 288
rect 348 252 360 288
rect 372 252 384 288
rect 396 285 408 288
rect 396 279 399 285
rect 405 279 408 285
rect 396 273 408 279
rect 396 267 399 273
rect 405 267 408 273
rect 396 261 408 267
rect 396 255 399 261
rect 405 255 408 261
rect 396 252 408 255
rect 420 285 432 288
rect 420 279 423 285
rect 429 279 432 285
rect 420 273 432 279
rect 420 267 423 273
rect 429 267 432 273
rect 420 261 432 267
rect 420 255 423 261
rect 429 255 432 261
rect 420 252 432 255
rect 444 252 456 288
rect 468 252 480 288
rect 492 252 504 288
rect 516 285 528 288
rect 516 279 519 285
rect 525 279 528 285
rect 516 273 528 279
rect 516 267 519 273
rect 525 267 528 273
rect 516 261 528 267
rect 516 255 519 261
rect 525 255 528 261
rect 516 252 528 255
rect 540 252 552 288
rect 564 252 576 288
rect 588 252 600 288
rect 612 285 624 288
rect 612 279 615 285
rect 621 279 624 285
rect 612 273 624 279
rect 612 267 615 273
rect 621 267 624 273
rect 612 261 624 267
rect 612 255 615 261
rect 621 255 624 261
rect 612 252 624 255
rect 636 285 648 288
rect 636 279 639 285
rect 645 279 648 285
rect 636 273 648 279
rect 636 267 639 273
rect 645 267 648 273
rect 636 261 648 267
rect 636 255 639 261
rect 645 255 648 261
rect 636 252 648 255
rect 660 252 672 288
rect 684 252 696 288
rect 708 252 720 288
rect 732 285 744 288
rect 732 279 735 285
rect 741 279 744 285
rect 732 273 744 279
rect 732 267 735 273
rect 741 267 744 273
rect 732 261 744 267
rect 732 255 735 261
rect 741 255 744 261
rect 732 252 744 255
rect 756 252 768 288
rect 780 252 792 288
rect 804 252 816 288
rect 828 285 840 288
rect 828 279 831 285
rect 837 279 840 285
rect 828 273 840 279
rect 828 267 831 273
rect 837 267 840 273
rect 828 261 840 267
rect 828 255 831 261
rect 837 255 840 261
rect 828 252 840 255
rect 852 285 864 288
rect 852 279 855 285
rect 861 279 864 285
rect 852 273 864 279
rect 852 267 855 273
rect 861 267 864 273
rect 852 261 864 267
rect 852 255 855 261
rect 861 255 864 261
rect 852 252 864 255
rect 876 285 888 288
rect 876 279 879 285
rect 885 279 888 285
rect 876 273 888 279
rect 876 267 879 273
rect 885 267 888 273
rect 876 261 888 267
rect 876 255 879 261
rect 885 255 888 261
rect 876 252 888 255
rect 900 285 912 288
rect 900 279 903 285
rect 909 279 912 285
rect 900 273 912 279
rect 900 267 903 273
rect 909 267 912 273
rect 900 261 912 267
rect 900 255 903 261
rect 909 255 912 261
rect 900 252 912 255
rect 924 252 936 288
rect 948 252 960 288
rect 972 252 984 288
rect 996 252 1008 288
rect 1020 252 1032 288
rect 1044 285 1056 288
rect 1044 279 1047 285
rect 1053 279 1056 285
rect 1044 273 1056 279
rect 1044 267 1047 273
rect 1053 267 1056 273
rect 1044 261 1056 267
rect 1044 255 1047 261
rect 1053 255 1056 261
rect 1044 252 1056 255
rect 1068 285 1080 288
rect 1068 279 1071 285
rect 1077 279 1080 285
rect 1068 273 1080 279
rect 1068 267 1071 273
rect 1077 267 1080 273
rect 1068 261 1080 267
rect 1068 255 1071 261
rect 1077 255 1080 261
rect 1068 252 1080 255
rect 1092 285 1104 288
rect 1092 279 1095 285
rect 1101 279 1104 285
rect 1092 273 1104 279
rect 1092 267 1095 273
rect 1101 267 1104 273
rect 1092 261 1104 267
rect 1092 255 1095 261
rect 1101 255 1104 261
rect 1092 252 1104 255
rect 1116 285 1128 288
rect 1116 279 1119 285
rect 1125 279 1128 285
rect 1116 273 1128 279
rect 1116 267 1119 273
rect 1125 267 1128 273
rect 1116 261 1128 267
rect 1116 255 1119 261
rect 1125 255 1128 261
rect 1116 252 1128 255
rect 1140 285 1152 288
rect 1140 279 1143 285
rect 1149 279 1152 285
rect 1140 273 1152 279
rect 1140 267 1143 273
rect 1149 267 1152 273
rect 1140 261 1152 267
rect 1140 255 1143 261
rect 1149 255 1152 261
rect 1140 252 1152 255
rect 1164 285 1176 288
rect 1164 279 1167 285
rect 1173 279 1176 285
rect 1164 273 1176 279
rect 1164 267 1167 273
rect 1173 267 1176 273
rect 1164 261 1176 267
rect 1164 255 1167 261
rect 1173 255 1176 261
rect 1164 252 1176 255
rect 1188 285 1200 288
rect 1188 279 1191 285
rect 1197 279 1200 285
rect 1188 273 1200 279
rect 1188 267 1191 273
rect 1197 267 1200 273
rect 1188 261 1200 267
rect 1188 255 1191 261
rect 1197 255 1200 261
rect 1188 252 1200 255
rect 1212 285 1224 288
rect 1212 279 1215 285
rect 1221 279 1224 285
rect 1212 273 1224 279
rect 1212 267 1215 273
rect 1221 267 1224 273
rect 1212 261 1224 267
rect 1212 255 1215 261
rect 1221 255 1224 261
rect 1212 252 1224 255
rect 1236 285 1248 288
rect 1236 279 1239 285
rect 1245 279 1248 285
rect 1236 273 1248 279
rect 1236 267 1239 273
rect 1245 267 1248 273
rect 1236 261 1248 267
rect 1236 255 1239 261
rect 1245 255 1248 261
rect 1236 252 1248 255
rect 1260 285 1272 288
rect 1260 279 1263 285
rect 1269 279 1272 285
rect 1260 273 1272 279
rect 1260 267 1263 273
rect 1269 267 1272 273
rect 1260 261 1272 267
rect 1260 255 1263 261
rect 1269 255 1272 261
rect 1260 252 1272 255
rect 1284 285 1296 288
rect 1284 279 1287 285
rect 1293 279 1296 285
rect 1284 273 1296 279
rect 1284 267 1287 273
rect 1293 267 1296 273
rect 1284 261 1296 267
rect 1284 255 1287 261
rect 1293 255 1296 261
rect 1284 252 1296 255
rect 1308 285 1320 288
rect 1308 279 1311 285
rect 1317 279 1320 285
rect 1308 273 1320 279
rect 1308 267 1311 273
rect 1317 267 1320 273
rect 1308 261 1320 267
rect 1308 255 1311 261
rect 1317 255 1320 261
rect 1308 252 1320 255
rect 1332 285 1344 288
rect 1332 279 1335 285
rect 1341 279 1344 285
rect 1332 273 1344 279
rect 1332 267 1335 273
rect 1341 267 1344 273
rect 1332 261 1344 267
rect 1332 255 1335 261
rect 1341 255 1344 261
rect 1332 252 1344 255
rect 1356 285 1368 288
rect 1356 279 1359 285
rect 1365 279 1368 285
rect 1356 273 1368 279
rect 1356 267 1359 273
rect 1365 267 1368 273
rect 1356 261 1368 267
rect 1356 255 1359 261
rect 1365 255 1368 261
rect 1356 252 1368 255
rect 1380 285 1392 288
rect 1380 279 1383 285
rect 1389 279 1392 285
rect 1380 273 1392 279
rect 1380 267 1383 273
rect 1389 267 1392 273
rect 1380 261 1392 267
rect 1380 255 1383 261
rect 1389 255 1392 261
rect 1380 252 1392 255
rect 1404 285 1416 288
rect 1404 279 1407 285
rect 1413 279 1416 285
rect 1404 273 1416 279
rect 1404 267 1407 273
rect 1413 267 1416 273
rect 1404 261 1416 267
rect 1404 255 1407 261
rect 1413 255 1416 261
rect 1404 252 1416 255
rect 1428 285 1440 288
rect 1428 279 1431 285
rect 1437 279 1440 285
rect 1428 273 1440 279
rect 1428 267 1431 273
rect 1437 267 1440 273
rect 1428 261 1440 267
rect 1428 255 1431 261
rect 1437 255 1440 261
rect 1428 252 1440 255
rect 1452 285 1464 288
rect 1452 279 1455 285
rect 1461 279 1464 285
rect 1452 273 1464 279
rect 1452 267 1455 273
rect 1461 267 1464 273
rect 1452 261 1464 267
rect 1452 255 1455 261
rect 1461 255 1464 261
rect 1452 252 1464 255
rect 1476 285 1488 288
rect 1476 279 1479 285
rect 1485 279 1488 285
rect 1476 273 1488 279
rect 1476 267 1479 273
rect 1485 267 1488 273
rect 1476 261 1488 267
rect 1476 255 1479 261
rect 1485 255 1488 261
rect 1476 252 1488 255
<< mvpdiff >>
rect -12 573 0 576
rect -12 567 -9 573
rect -3 567 0 573
rect -12 561 0 567
rect -12 555 -9 561
rect -3 555 0 561
rect -12 549 0 555
rect -12 543 -9 549
rect -3 543 0 549
rect -12 540 0 543
rect 12 573 24 576
rect 12 567 15 573
rect 21 567 24 573
rect 12 561 24 567
rect 12 555 15 561
rect 21 555 24 561
rect 12 549 24 555
rect 12 543 15 549
rect 21 543 24 549
rect 12 540 24 543
rect 36 573 48 576
rect 36 567 39 573
rect 45 567 48 573
rect 36 561 48 567
rect 36 555 39 561
rect 45 555 48 561
rect 36 549 48 555
rect 36 543 39 549
rect 45 543 48 549
rect 36 540 48 543
rect 60 573 72 576
rect 60 567 63 573
rect 69 567 72 573
rect 60 561 72 567
rect 60 555 63 561
rect 69 555 72 561
rect 60 549 72 555
rect 60 543 63 549
rect 69 543 72 549
rect 60 540 72 543
rect 84 573 96 576
rect 84 567 87 573
rect 93 567 96 573
rect 84 561 96 567
rect 84 555 87 561
rect 93 555 96 561
rect 84 549 96 555
rect 84 543 87 549
rect 93 543 96 549
rect 84 540 96 543
rect 108 573 120 576
rect 108 567 111 573
rect 117 567 120 573
rect 108 561 120 567
rect 108 555 111 561
rect 117 555 120 561
rect 108 549 120 555
rect 108 543 111 549
rect 117 543 120 549
rect 108 540 120 543
rect 132 573 144 576
rect 132 567 135 573
rect 141 567 144 573
rect 132 561 144 567
rect 132 555 135 561
rect 141 555 144 561
rect 132 549 144 555
rect 132 543 135 549
rect 141 543 144 549
rect 132 540 144 543
rect 156 573 168 576
rect 156 567 159 573
rect 165 567 168 573
rect 156 561 168 567
rect 156 555 159 561
rect 165 555 168 561
rect 156 549 168 555
rect 156 543 159 549
rect 165 543 168 549
rect 156 540 168 543
rect 180 573 192 576
rect 180 567 183 573
rect 189 567 192 573
rect 180 561 192 567
rect 180 555 183 561
rect 189 555 192 561
rect 180 549 192 555
rect 180 543 183 549
rect 189 543 192 549
rect 180 540 192 543
rect 204 573 216 576
rect 204 567 207 573
rect 213 567 216 573
rect 204 561 216 567
rect 204 555 207 561
rect 213 555 216 561
rect 204 549 216 555
rect 204 543 207 549
rect 213 543 216 549
rect 204 540 216 543
rect 228 540 240 576
rect 252 573 264 576
rect 252 567 255 573
rect 261 567 264 573
rect 252 561 264 567
rect 252 555 255 561
rect 261 555 264 561
rect 252 549 264 555
rect 252 543 255 549
rect 261 543 264 549
rect 252 540 264 543
rect 276 540 288 576
rect 300 573 312 576
rect 300 567 303 573
rect 309 567 312 573
rect 300 561 312 567
rect 300 555 303 561
rect 309 555 312 561
rect 300 549 312 555
rect 300 543 303 549
rect 309 543 312 549
rect 300 540 312 543
rect 324 540 336 576
rect 348 573 360 576
rect 348 567 351 573
rect 357 567 360 573
rect 348 561 360 567
rect 348 555 351 561
rect 357 555 360 561
rect 348 549 360 555
rect 348 543 351 549
rect 357 543 360 549
rect 348 540 360 543
rect 372 540 384 576
rect 396 573 408 576
rect 396 567 399 573
rect 405 567 408 573
rect 396 561 408 567
rect 396 555 399 561
rect 405 555 408 561
rect 396 549 408 555
rect 396 543 399 549
rect 405 543 408 549
rect 396 540 408 543
rect 420 573 432 576
rect 420 567 423 573
rect 429 567 432 573
rect 420 561 432 567
rect 420 555 423 561
rect 429 555 432 561
rect 420 549 432 555
rect 420 543 423 549
rect 429 543 432 549
rect 420 540 432 543
rect 444 540 456 576
rect 468 573 480 576
rect 468 567 471 573
rect 477 567 480 573
rect 468 561 480 567
rect 468 555 471 561
rect 477 555 480 561
rect 468 549 480 555
rect 468 543 471 549
rect 477 543 480 549
rect 468 540 480 543
rect 492 540 504 576
rect 516 573 528 576
rect 516 567 519 573
rect 525 567 528 573
rect 516 561 528 567
rect 516 555 519 561
rect 525 555 528 561
rect 516 549 528 555
rect 516 543 519 549
rect 525 543 528 549
rect 516 540 528 543
rect 540 540 552 576
rect 564 573 576 576
rect 564 567 567 573
rect 573 567 576 573
rect 564 561 576 567
rect 564 555 567 561
rect 573 555 576 561
rect 564 549 576 555
rect 564 543 567 549
rect 573 543 576 549
rect 564 540 576 543
rect 588 540 600 576
rect 612 573 624 576
rect 612 567 615 573
rect 621 567 624 573
rect 612 561 624 567
rect 612 555 615 561
rect 621 555 624 561
rect 612 549 624 555
rect 612 543 615 549
rect 621 543 624 549
rect 612 540 624 543
rect 636 573 648 576
rect 636 567 639 573
rect 645 567 648 573
rect 636 561 648 567
rect 636 555 639 561
rect 645 555 648 561
rect 636 549 648 555
rect 636 543 639 549
rect 645 543 648 549
rect 636 540 648 543
rect 660 540 672 576
rect 684 540 696 576
rect 708 540 720 576
rect 732 540 744 576
rect 756 540 768 576
rect 780 540 792 576
rect 804 540 816 576
rect 828 573 840 576
rect 828 567 831 573
rect 837 567 840 573
rect 828 561 840 567
rect 828 555 831 561
rect 837 555 840 561
rect 828 549 840 555
rect 828 543 831 549
rect 837 543 840 549
rect 828 540 840 543
rect 852 573 864 576
rect 852 567 855 573
rect 861 567 864 573
rect 852 561 864 567
rect 852 555 855 561
rect 861 555 864 561
rect 852 549 864 555
rect 852 543 855 549
rect 861 543 864 549
rect 852 540 864 543
rect 876 540 888 576
rect 900 540 912 576
rect 924 540 936 576
rect 948 540 960 576
rect 972 540 984 576
rect 996 540 1008 576
rect 1020 540 1032 576
rect 1044 573 1056 576
rect 1044 567 1047 573
rect 1053 567 1056 573
rect 1044 561 1056 567
rect 1044 555 1047 561
rect 1053 555 1056 561
rect 1044 549 1056 555
rect 1044 543 1047 549
rect 1053 543 1056 549
rect 1044 540 1056 543
rect 1068 573 1080 576
rect 1068 567 1071 573
rect 1077 567 1080 573
rect 1068 561 1080 567
rect 1068 555 1071 561
rect 1077 555 1080 561
rect 1068 549 1080 555
rect 1068 543 1071 549
rect 1077 543 1080 549
rect 1068 540 1080 543
rect 1092 573 1104 576
rect 1092 567 1095 573
rect 1101 567 1104 573
rect 1092 561 1104 567
rect 1092 555 1095 561
rect 1101 555 1104 561
rect 1092 549 1104 555
rect 1092 543 1095 549
rect 1101 543 1104 549
rect 1092 540 1104 543
rect 1116 573 1128 576
rect 1116 567 1119 573
rect 1125 567 1128 573
rect 1116 561 1128 567
rect 1116 555 1119 561
rect 1125 555 1128 561
rect 1116 549 1128 555
rect 1116 543 1119 549
rect 1125 543 1128 549
rect 1116 540 1128 543
rect 1140 573 1152 576
rect 1140 567 1143 573
rect 1149 567 1152 573
rect 1140 561 1152 567
rect 1140 555 1143 561
rect 1149 555 1152 561
rect 1140 549 1152 555
rect 1140 543 1143 549
rect 1149 543 1152 549
rect 1140 540 1152 543
rect 1164 573 1176 576
rect 1164 567 1167 573
rect 1173 567 1176 573
rect 1164 561 1176 567
rect 1164 555 1167 561
rect 1173 555 1176 561
rect 1164 549 1176 555
rect 1164 543 1167 549
rect 1173 543 1176 549
rect 1164 540 1176 543
rect 1188 573 1200 576
rect 1188 567 1191 573
rect 1197 567 1200 573
rect 1188 561 1200 567
rect 1188 555 1191 561
rect 1197 555 1200 561
rect 1188 549 1200 555
rect 1188 543 1191 549
rect 1197 543 1200 549
rect 1188 540 1200 543
rect 1212 573 1224 576
rect 1212 567 1215 573
rect 1221 567 1224 573
rect 1212 561 1224 567
rect 1212 555 1215 561
rect 1221 555 1224 561
rect 1212 549 1224 555
rect 1212 543 1215 549
rect 1221 543 1224 549
rect 1212 540 1224 543
rect 1236 573 1248 576
rect 1236 567 1239 573
rect 1245 567 1248 573
rect 1236 561 1248 567
rect 1236 555 1239 561
rect 1245 555 1248 561
rect 1236 549 1248 555
rect 1236 543 1239 549
rect 1245 543 1248 549
rect 1236 540 1248 543
rect 1260 573 1272 576
rect 1260 567 1263 573
rect 1269 567 1272 573
rect 1260 561 1272 567
rect 1260 555 1263 561
rect 1269 555 1272 561
rect 1260 549 1272 555
rect 1260 543 1263 549
rect 1269 543 1272 549
rect 1260 540 1272 543
rect 1284 573 1296 576
rect 1284 567 1287 573
rect 1293 567 1296 573
rect 1284 561 1296 567
rect 1284 555 1287 561
rect 1293 555 1296 561
rect 1284 549 1296 555
rect 1284 543 1287 549
rect 1293 543 1296 549
rect 1284 540 1296 543
rect 1308 573 1320 576
rect 1308 567 1311 573
rect 1317 567 1320 573
rect 1308 561 1320 567
rect 1308 555 1311 561
rect 1317 555 1320 561
rect 1308 549 1320 555
rect 1308 543 1311 549
rect 1317 543 1320 549
rect 1308 540 1320 543
rect 1332 573 1344 576
rect 1332 567 1335 573
rect 1341 567 1344 573
rect 1332 561 1344 567
rect 1332 555 1335 561
rect 1341 555 1344 561
rect 1332 549 1344 555
rect 1332 543 1335 549
rect 1341 543 1344 549
rect 1332 540 1344 543
rect 1356 573 1368 576
rect 1356 567 1359 573
rect 1365 567 1368 573
rect 1356 561 1368 567
rect 1356 555 1359 561
rect 1365 555 1368 561
rect 1356 549 1368 555
rect 1356 543 1359 549
rect 1365 543 1368 549
rect 1356 540 1368 543
rect 1380 573 1392 576
rect 1380 567 1383 573
rect 1389 567 1392 573
rect 1380 561 1392 567
rect 1380 555 1383 561
rect 1389 555 1392 561
rect 1380 549 1392 555
rect 1380 543 1383 549
rect 1389 543 1392 549
rect 1380 540 1392 543
rect 1404 573 1416 576
rect 1404 567 1407 573
rect 1413 567 1416 573
rect 1404 561 1416 567
rect 1404 555 1407 561
rect 1413 555 1416 561
rect 1404 549 1416 555
rect 1404 543 1407 549
rect 1413 543 1416 549
rect 1404 540 1416 543
rect 1428 573 1440 576
rect 1428 567 1431 573
rect 1437 567 1440 573
rect 1428 561 1440 567
rect 1428 555 1431 561
rect 1437 555 1440 561
rect 1428 549 1440 555
rect 1428 543 1431 549
rect 1437 543 1440 549
rect 1428 540 1440 543
rect 1452 573 1464 576
rect 1452 567 1455 573
rect 1461 567 1464 573
rect 1452 561 1464 567
rect 1452 555 1455 561
rect 1461 555 1464 561
rect 1452 549 1464 555
rect 1452 543 1455 549
rect 1461 543 1464 549
rect 1452 540 1464 543
rect 1476 573 1488 576
rect 1476 567 1479 573
rect 1485 567 1488 573
rect 1476 561 1488 567
rect 1476 555 1479 561
rect 1485 555 1488 561
rect 1476 549 1488 555
rect 1476 543 1479 549
rect 1485 543 1488 549
rect 1476 540 1488 543
rect -12 477 0 480
rect -12 471 -9 477
rect -3 471 0 477
rect -12 465 0 471
rect -12 459 -9 465
rect -3 459 0 465
rect -12 453 0 459
rect -12 447 -9 453
rect -3 447 0 453
rect -12 444 0 447
rect 12 477 24 480
rect 12 471 15 477
rect 21 471 24 477
rect 12 465 24 471
rect 12 459 15 465
rect 21 459 24 465
rect 12 453 24 459
rect 12 447 15 453
rect 21 447 24 453
rect 12 444 24 447
rect 36 477 48 480
rect 36 471 39 477
rect 45 471 48 477
rect 36 465 48 471
rect 36 459 39 465
rect 45 459 48 465
rect 36 453 48 459
rect 36 447 39 453
rect 45 447 48 453
rect 36 444 48 447
rect 60 477 72 480
rect 60 471 63 477
rect 69 471 72 477
rect 60 465 72 471
rect 60 459 63 465
rect 69 459 72 465
rect 60 453 72 459
rect 60 447 63 453
rect 69 447 72 453
rect 60 444 72 447
rect 84 477 96 480
rect 84 471 87 477
rect 93 471 96 477
rect 84 465 96 471
rect 84 459 87 465
rect 93 459 96 465
rect 84 453 96 459
rect 84 447 87 453
rect 93 447 96 453
rect 84 444 96 447
rect 108 477 120 480
rect 108 471 111 477
rect 117 471 120 477
rect 108 465 120 471
rect 108 459 111 465
rect 117 459 120 465
rect 108 453 120 459
rect 108 447 111 453
rect 117 447 120 453
rect 108 444 120 447
rect 132 477 144 480
rect 132 471 135 477
rect 141 471 144 477
rect 132 465 144 471
rect 132 459 135 465
rect 141 459 144 465
rect 132 453 144 459
rect 132 447 135 453
rect 141 447 144 453
rect 132 444 144 447
rect 156 477 168 480
rect 156 471 159 477
rect 165 471 168 477
rect 156 465 168 471
rect 156 459 159 465
rect 165 459 168 465
rect 156 453 168 459
rect 156 447 159 453
rect 165 447 168 453
rect 156 444 168 447
rect 180 477 192 480
rect 180 471 183 477
rect 189 471 192 477
rect 180 465 192 471
rect 180 459 183 465
rect 189 459 192 465
rect 180 453 192 459
rect 180 447 183 453
rect 189 447 192 453
rect 180 444 192 447
rect 204 477 216 480
rect 204 471 207 477
rect 213 471 216 477
rect 204 465 216 471
rect 204 459 207 465
rect 213 459 216 465
rect 204 453 216 459
rect 204 447 207 453
rect 213 447 216 453
rect 204 444 216 447
rect 228 444 240 480
rect 252 477 264 480
rect 252 471 255 477
rect 261 471 264 477
rect 252 465 264 471
rect 252 459 255 465
rect 261 459 264 465
rect 252 453 264 459
rect 252 447 255 453
rect 261 447 264 453
rect 252 444 264 447
rect 276 444 288 480
rect 300 477 312 480
rect 300 471 303 477
rect 309 471 312 477
rect 300 465 312 471
rect 300 459 303 465
rect 309 459 312 465
rect 300 453 312 459
rect 300 447 303 453
rect 309 447 312 453
rect 300 444 312 447
rect 324 444 336 480
rect 348 477 360 480
rect 348 471 351 477
rect 357 471 360 477
rect 348 465 360 471
rect 348 459 351 465
rect 357 459 360 465
rect 348 453 360 459
rect 348 447 351 453
rect 357 447 360 453
rect 348 444 360 447
rect 372 444 384 480
rect 396 477 408 480
rect 396 471 399 477
rect 405 471 408 477
rect 396 465 408 471
rect 396 459 399 465
rect 405 459 408 465
rect 396 453 408 459
rect 396 447 399 453
rect 405 447 408 453
rect 396 444 408 447
rect 420 477 432 480
rect 420 471 423 477
rect 429 471 432 477
rect 420 465 432 471
rect 420 459 423 465
rect 429 459 432 465
rect 420 453 432 459
rect 420 447 423 453
rect 429 447 432 453
rect 420 444 432 447
rect 444 444 456 480
rect 468 477 480 480
rect 468 471 471 477
rect 477 471 480 477
rect 468 465 480 471
rect 468 459 471 465
rect 477 459 480 465
rect 468 453 480 459
rect 468 447 471 453
rect 477 447 480 453
rect 468 444 480 447
rect 492 444 504 480
rect 516 477 528 480
rect 516 471 519 477
rect 525 471 528 477
rect 516 465 528 471
rect 516 459 519 465
rect 525 459 528 465
rect 516 453 528 459
rect 516 447 519 453
rect 525 447 528 453
rect 516 444 528 447
rect 540 444 552 480
rect 564 477 576 480
rect 564 471 567 477
rect 573 471 576 477
rect 564 465 576 471
rect 564 459 567 465
rect 573 459 576 465
rect 564 453 576 459
rect 564 447 567 453
rect 573 447 576 453
rect 564 444 576 447
rect 588 444 600 480
rect 612 477 624 480
rect 612 471 615 477
rect 621 471 624 477
rect 612 465 624 471
rect 612 459 615 465
rect 621 459 624 465
rect 612 453 624 459
rect 612 447 615 453
rect 621 447 624 453
rect 612 444 624 447
rect 636 477 648 480
rect 636 471 639 477
rect 645 471 648 477
rect 636 465 648 471
rect 636 459 639 465
rect 645 459 648 465
rect 636 453 648 459
rect 636 447 639 453
rect 645 447 648 453
rect 636 444 648 447
rect 660 444 672 480
rect 684 444 696 480
rect 708 444 720 480
rect 732 444 744 480
rect 756 444 768 480
rect 780 444 792 480
rect 804 444 816 480
rect 828 477 840 480
rect 828 471 831 477
rect 837 471 840 477
rect 828 465 840 471
rect 828 459 831 465
rect 837 459 840 465
rect 828 453 840 459
rect 828 447 831 453
rect 837 447 840 453
rect 828 444 840 447
rect 852 477 864 480
rect 852 471 855 477
rect 861 471 864 477
rect 852 465 864 471
rect 852 459 855 465
rect 861 459 864 465
rect 852 453 864 459
rect 852 447 855 453
rect 861 447 864 453
rect 852 444 864 447
rect 876 444 888 480
rect 900 444 912 480
rect 924 444 936 480
rect 948 444 960 480
rect 972 444 984 480
rect 996 444 1008 480
rect 1020 444 1032 480
rect 1044 477 1056 480
rect 1044 471 1047 477
rect 1053 471 1056 477
rect 1044 465 1056 471
rect 1044 459 1047 465
rect 1053 459 1056 465
rect 1044 453 1056 459
rect 1044 447 1047 453
rect 1053 447 1056 453
rect 1044 444 1056 447
rect 1068 477 1080 480
rect 1068 471 1071 477
rect 1077 471 1080 477
rect 1068 465 1080 471
rect 1068 459 1071 465
rect 1077 459 1080 465
rect 1068 453 1080 459
rect 1068 447 1071 453
rect 1077 447 1080 453
rect 1068 444 1080 447
rect 1092 477 1104 480
rect 1092 471 1095 477
rect 1101 471 1104 477
rect 1092 465 1104 471
rect 1092 459 1095 465
rect 1101 459 1104 465
rect 1092 453 1104 459
rect 1092 447 1095 453
rect 1101 447 1104 453
rect 1092 444 1104 447
rect 1116 477 1128 480
rect 1116 471 1119 477
rect 1125 471 1128 477
rect 1116 465 1128 471
rect 1116 459 1119 465
rect 1125 459 1128 465
rect 1116 453 1128 459
rect 1116 447 1119 453
rect 1125 447 1128 453
rect 1116 444 1128 447
rect 1140 477 1152 480
rect 1140 471 1143 477
rect 1149 471 1152 477
rect 1140 465 1152 471
rect 1140 459 1143 465
rect 1149 459 1152 465
rect 1140 453 1152 459
rect 1140 447 1143 453
rect 1149 447 1152 453
rect 1140 444 1152 447
rect 1164 477 1176 480
rect 1164 471 1167 477
rect 1173 471 1176 477
rect 1164 465 1176 471
rect 1164 459 1167 465
rect 1173 459 1176 465
rect 1164 453 1176 459
rect 1164 447 1167 453
rect 1173 447 1176 453
rect 1164 444 1176 447
rect 1188 477 1200 480
rect 1188 471 1191 477
rect 1197 471 1200 477
rect 1188 465 1200 471
rect 1188 459 1191 465
rect 1197 459 1200 465
rect 1188 453 1200 459
rect 1188 447 1191 453
rect 1197 447 1200 453
rect 1188 444 1200 447
rect 1212 477 1224 480
rect 1212 471 1215 477
rect 1221 471 1224 477
rect 1212 465 1224 471
rect 1212 459 1215 465
rect 1221 459 1224 465
rect 1212 453 1224 459
rect 1212 447 1215 453
rect 1221 447 1224 453
rect 1212 444 1224 447
rect 1236 477 1248 480
rect 1236 471 1239 477
rect 1245 471 1248 477
rect 1236 465 1248 471
rect 1236 459 1239 465
rect 1245 459 1248 465
rect 1236 453 1248 459
rect 1236 447 1239 453
rect 1245 447 1248 453
rect 1236 444 1248 447
rect 1260 477 1272 480
rect 1260 471 1263 477
rect 1269 471 1272 477
rect 1260 465 1272 471
rect 1260 459 1263 465
rect 1269 459 1272 465
rect 1260 453 1272 459
rect 1260 447 1263 453
rect 1269 447 1272 453
rect 1260 444 1272 447
rect 1284 477 1296 480
rect 1284 471 1287 477
rect 1293 471 1296 477
rect 1284 465 1296 471
rect 1284 459 1287 465
rect 1293 459 1296 465
rect 1284 453 1296 459
rect 1284 447 1287 453
rect 1293 447 1296 453
rect 1284 444 1296 447
rect 1308 477 1320 480
rect 1308 471 1311 477
rect 1317 471 1320 477
rect 1308 465 1320 471
rect 1308 459 1311 465
rect 1317 459 1320 465
rect 1308 453 1320 459
rect 1308 447 1311 453
rect 1317 447 1320 453
rect 1308 444 1320 447
rect 1332 477 1344 480
rect 1332 471 1335 477
rect 1341 471 1344 477
rect 1332 465 1344 471
rect 1332 459 1335 465
rect 1341 459 1344 465
rect 1332 453 1344 459
rect 1332 447 1335 453
rect 1341 447 1344 453
rect 1332 444 1344 447
rect 1356 477 1368 480
rect 1356 471 1359 477
rect 1365 471 1368 477
rect 1356 465 1368 471
rect 1356 459 1359 465
rect 1365 459 1368 465
rect 1356 453 1368 459
rect 1356 447 1359 453
rect 1365 447 1368 453
rect 1356 444 1368 447
rect 1380 477 1392 480
rect 1380 471 1383 477
rect 1389 471 1392 477
rect 1380 465 1392 471
rect 1380 459 1383 465
rect 1389 459 1392 465
rect 1380 453 1392 459
rect 1380 447 1383 453
rect 1389 447 1392 453
rect 1380 444 1392 447
rect 1404 477 1416 480
rect 1404 471 1407 477
rect 1413 471 1416 477
rect 1404 465 1416 471
rect 1404 459 1407 465
rect 1413 459 1416 465
rect 1404 453 1416 459
rect 1404 447 1407 453
rect 1413 447 1416 453
rect 1404 444 1416 447
rect 1428 477 1440 480
rect 1428 471 1431 477
rect 1437 471 1440 477
rect 1428 465 1440 471
rect 1428 459 1431 465
rect 1437 459 1440 465
rect 1428 453 1440 459
rect 1428 447 1431 453
rect 1437 447 1440 453
rect 1428 444 1440 447
rect 1452 477 1464 480
rect 1452 471 1455 477
rect 1461 471 1464 477
rect 1452 465 1464 471
rect 1452 459 1455 465
rect 1461 459 1464 465
rect 1452 453 1464 459
rect 1452 447 1455 453
rect 1461 447 1464 453
rect 1452 444 1464 447
rect 1476 477 1488 480
rect 1476 471 1479 477
rect 1485 471 1488 477
rect 1476 465 1488 471
rect 1476 459 1479 465
rect 1485 459 1488 465
rect 1476 453 1488 459
rect 1476 447 1479 453
rect 1485 447 1488 453
rect 1476 444 1488 447
<< ndiffc >>
rect -9 39 -3 45
rect -9 27 -3 33
rect -9 15 -3 21
rect 39 39 45 45
rect 39 27 45 33
rect 39 15 45 21
rect 87 39 93 45
rect 87 27 93 33
rect 87 15 93 21
rect 135 39 141 45
rect 135 27 141 33
rect 135 15 141 21
rect 183 39 189 45
rect 183 27 189 33
rect 183 15 189 21
rect 207 39 213 45
rect 207 27 213 33
rect 207 15 213 21
rect 255 39 261 45
rect 255 27 261 33
rect 255 15 261 21
rect 303 39 309 45
rect 303 27 309 33
rect 303 15 309 21
rect 351 39 357 45
rect 351 27 357 33
rect 351 15 357 21
rect 399 39 405 45
rect 399 27 405 33
rect 399 15 405 21
rect 423 39 429 45
rect 423 27 429 33
rect 423 15 429 21
rect 519 39 525 45
rect 519 27 525 33
rect 519 15 525 21
rect 615 39 621 45
rect 615 27 621 33
rect 615 15 621 21
rect 639 39 645 45
rect 639 27 645 33
rect 639 15 645 21
rect 735 39 741 45
rect 735 27 741 33
rect 735 15 741 21
rect 831 39 837 45
rect 831 27 837 33
rect 831 15 837 21
rect 855 39 861 45
rect 855 27 861 33
rect 855 15 861 21
rect 1047 39 1053 45
rect 1047 27 1053 33
rect 1047 15 1053 21
rect 1071 39 1077 45
rect 1071 27 1077 33
rect 1071 15 1077 21
rect 1095 39 1101 45
rect 1095 27 1101 33
rect 1095 15 1101 21
rect 1119 39 1125 45
rect 1119 27 1125 33
rect 1119 15 1125 21
rect 1143 39 1149 45
rect 1143 27 1149 33
rect 1143 15 1149 21
rect 1167 39 1173 45
rect 1167 27 1173 33
rect 1167 15 1173 21
rect 1191 39 1197 45
rect 1191 27 1197 33
rect 1191 15 1197 21
rect 1215 39 1221 45
rect 1215 27 1221 33
rect 1215 15 1221 21
rect 1239 39 1245 45
rect 1239 27 1245 33
rect 1239 15 1245 21
rect 1263 39 1269 45
rect 1263 27 1269 33
rect 1263 15 1269 21
rect 1287 39 1293 45
rect 1287 27 1293 33
rect 1287 15 1293 21
rect 1311 39 1317 45
rect 1311 27 1317 33
rect 1311 15 1317 21
rect 1335 39 1341 45
rect 1335 27 1341 33
rect 1335 15 1341 21
rect 1359 39 1365 45
rect 1359 27 1365 33
rect 1359 15 1365 21
rect 1383 39 1389 45
rect 1383 27 1389 33
rect 1383 15 1389 21
rect 1407 39 1413 45
rect 1407 27 1413 33
rect 1407 15 1413 21
rect 1431 39 1437 45
rect 1431 27 1437 33
rect 1431 15 1437 21
rect 1455 39 1461 45
rect 1455 27 1461 33
rect 1455 15 1461 21
rect 1479 39 1485 45
rect 1479 27 1485 33
rect 1479 15 1485 21
<< mvndiffc >>
rect -9 279 -3 285
rect -9 267 -3 273
rect -9 255 -3 261
rect 15 279 21 285
rect 15 267 21 273
rect 15 255 21 261
rect 39 279 45 285
rect 39 267 45 273
rect 39 255 45 261
rect 63 279 69 285
rect 63 267 69 273
rect 63 255 69 261
rect 87 279 93 285
rect 87 267 93 273
rect 87 255 93 261
rect 111 279 117 285
rect 111 267 117 273
rect 111 255 117 261
rect 135 279 141 285
rect 135 267 141 273
rect 135 255 141 261
rect 159 279 165 285
rect 159 267 165 273
rect 159 255 165 261
rect 183 279 189 285
rect 183 267 189 273
rect 183 255 189 261
rect 207 279 213 285
rect 207 267 213 273
rect 207 255 213 261
rect 303 279 309 285
rect 303 267 309 273
rect 303 255 309 261
rect 399 279 405 285
rect 399 267 405 273
rect 399 255 405 261
rect 423 279 429 285
rect 423 267 429 273
rect 423 255 429 261
rect 519 279 525 285
rect 519 267 525 273
rect 519 255 525 261
rect 615 279 621 285
rect 615 267 621 273
rect 615 255 621 261
rect 639 279 645 285
rect 639 267 645 273
rect 639 255 645 261
rect 735 279 741 285
rect 735 267 741 273
rect 735 255 741 261
rect 831 279 837 285
rect 831 267 837 273
rect 831 255 837 261
rect 855 279 861 285
rect 855 267 861 273
rect 855 255 861 261
rect 879 279 885 285
rect 879 267 885 273
rect 879 255 885 261
rect 903 279 909 285
rect 903 267 909 273
rect 903 255 909 261
rect 1047 279 1053 285
rect 1047 267 1053 273
rect 1047 255 1053 261
rect 1071 279 1077 285
rect 1071 267 1077 273
rect 1071 255 1077 261
rect 1095 279 1101 285
rect 1095 267 1101 273
rect 1095 255 1101 261
rect 1119 279 1125 285
rect 1119 267 1125 273
rect 1119 255 1125 261
rect 1143 279 1149 285
rect 1143 267 1149 273
rect 1143 255 1149 261
rect 1167 279 1173 285
rect 1167 267 1173 273
rect 1167 255 1173 261
rect 1191 279 1197 285
rect 1191 267 1197 273
rect 1191 255 1197 261
rect 1215 279 1221 285
rect 1215 267 1221 273
rect 1215 255 1221 261
rect 1239 279 1245 285
rect 1239 267 1245 273
rect 1239 255 1245 261
rect 1263 279 1269 285
rect 1263 267 1269 273
rect 1263 255 1269 261
rect 1287 279 1293 285
rect 1287 267 1293 273
rect 1287 255 1293 261
rect 1311 279 1317 285
rect 1311 267 1317 273
rect 1311 255 1317 261
rect 1335 279 1341 285
rect 1335 267 1341 273
rect 1335 255 1341 261
rect 1359 279 1365 285
rect 1359 267 1365 273
rect 1359 255 1365 261
rect 1383 279 1389 285
rect 1383 267 1389 273
rect 1383 255 1389 261
rect 1407 279 1413 285
rect 1407 267 1413 273
rect 1407 255 1413 261
rect 1431 279 1437 285
rect 1431 267 1437 273
rect 1431 255 1437 261
rect 1455 279 1461 285
rect 1455 267 1461 273
rect 1455 255 1461 261
rect 1479 279 1485 285
rect 1479 267 1485 273
rect 1479 255 1485 261
<< mvpdiffc >>
rect -9 567 -3 573
rect -9 555 -3 561
rect -9 543 -3 549
rect 15 567 21 573
rect 15 555 21 561
rect 15 543 21 549
rect 39 567 45 573
rect 39 555 45 561
rect 39 543 45 549
rect 63 567 69 573
rect 63 555 69 561
rect 63 543 69 549
rect 87 567 93 573
rect 87 555 93 561
rect 87 543 93 549
rect 111 567 117 573
rect 111 555 117 561
rect 111 543 117 549
rect 135 567 141 573
rect 135 555 141 561
rect 135 543 141 549
rect 159 567 165 573
rect 159 555 165 561
rect 159 543 165 549
rect 183 567 189 573
rect 183 555 189 561
rect 183 543 189 549
rect 207 567 213 573
rect 207 555 213 561
rect 207 543 213 549
rect 255 567 261 573
rect 255 555 261 561
rect 255 543 261 549
rect 303 567 309 573
rect 303 555 309 561
rect 303 543 309 549
rect 351 567 357 573
rect 351 555 357 561
rect 351 543 357 549
rect 399 567 405 573
rect 399 555 405 561
rect 399 543 405 549
rect 423 567 429 573
rect 423 555 429 561
rect 423 543 429 549
rect 471 567 477 573
rect 471 555 477 561
rect 471 543 477 549
rect 519 567 525 573
rect 519 555 525 561
rect 519 543 525 549
rect 567 567 573 573
rect 567 555 573 561
rect 567 543 573 549
rect 615 567 621 573
rect 615 555 621 561
rect 615 543 621 549
rect 639 567 645 573
rect 639 555 645 561
rect 639 543 645 549
rect 831 567 837 573
rect 831 555 837 561
rect 831 543 837 549
rect 855 567 861 573
rect 855 555 861 561
rect 855 543 861 549
rect 1047 567 1053 573
rect 1047 555 1053 561
rect 1047 543 1053 549
rect 1071 567 1077 573
rect 1071 555 1077 561
rect 1071 543 1077 549
rect 1095 567 1101 573
rect 1095 555 1101 561
rect 1095 543 1101 549
rect 1119 567 1125 573
rect 1119 555 1125 561
rect 1119 543 1125 549
rect 1143 567 1149 573
rect 1143 555 1149 561
rect 1143 543 1149 549
rect 1167 567 1173 573
rect 1167 555 1173 561
rect 1167 543 1173 549
rect 1191 567 1197 573
rect 1191 555 1197 561
rect 1191 543 1197 549
rect 1215 567 1221 573
rect 1215 555 1221 561
rect 1215 543 1221 549
rect 1239 567 1245 573
rect 1239 555 1245 561
rect 1239 543 1245 549
rect 1263 567 1269 573
rect 1263 555 1269 561
rect 1263 543 1269 549
rect 1287 567 1293 573
rect 1287 555 1293 561
rect 1287 543 1293 549
rect 1311 567 1317 573
rect 1311 555 1317 561
rect 1311 543 1317 549
rect 1335 567 1341 573
rect 1335 555 1341 561
rect 1335 543 1341 549
rect 1359 567 1365 573
rect 1359 555 1365 561
rect 1359 543 1365 549
rect 1383 567 1389 573
rect 1383 555 1389 561
rect 1383 543 1389 549
rect 1407 567 1413 573
rect 1407 555 1413 561
rect 1407 543 1413 549
rect 1431 567 1437 573
rect 1431 555 1437 561
rect 1431 543 1437 549
rect 1455 567 1461 573
rect 1455 555 1461 561
rect 1455 543 1461 549
rect 1479 567 1485 573
rect 1479 555 1485 561
rect 1479 543 1485 549
rect -9 471 -3 477
rect -9 459 -3 465
rect -9 447 -3 453
rect 15 471 21 477
rect 15 459 21 465
rect 15 447 21 453
rect 39 471 45 477
rect 39 459 45 465
rect 39 447 45 453
rect 63 471 69 477
rect 63 459 69 465
rect 63 447 69 453
rect 87 471 93 477
rect 87 459 93 465
rect 87 447 93 453
rect 111 471 117 477
rect 111 459 117 465
rect 111 447 117 453
rect 135 471 141 477
rect 135 459 141 465
rect 135 447 141 453
rect 159 471 165 477
rect 159 459 165 465
rect 159 447 165 453
rect 183 471 189 477
rect 183 459 189 465
rect 183 447 189 453
rect 207 471 213 477
rect 207 459 213 465
rect 207 447 213 453
rect 255 471 261 477
rect 255 459 261 465
rect 255 447 261 453
rect 303 471 309 477
rect 303 459 309 465
rect 303 447 309 453
rect 351 471 357 477
rect 351 459 357 465
rect 351 447 357 453
rect 399 471 405 477
rect 399 459 405 465
rect 399 447 405 453
rect 423 471 429 477
rect 423 459 429 465
rect 423 447 429 453
rect 471 471 477 477
rect 471 459 477 465
rect 471 447 477 453
rect 519 471 525 477
rect 519 459 525 465
rect 519 447 525 453
rect 567 471 573 477
rect 567 459 573 465
rect 567 447 573 453
rect 615 471 621 477
rect 615 459 621 465
rect 615 447 621 453
rect 639 471 645 477
rect 639 459 645 465
rect 639 447 645 453
rect 831 471 837 477
rect 831 459 837 465
rect 831 447 837 453
rect 855 471 861 477
rect 855 459 861 465
rect 855 447 861 453
rect 1047 471 1053 477
rect 1047 459 1053 465
rect 1047 447 1053 453
rect 1071 471 1077 477
rect 1071 459 1077 465
rect 1071 447 1077 453
rect 1095 471 1101 477
rect 1095 459 1101 465
rect 1095 447 1101 453
rect 1119 471 1125 477
rect 1119 459 1125 465
rect 1119 447 1125 453
rect 1143 471 1149 477
rect 1143 459 1149 465
rect 1143 447 1149 453
rect 1167 471 1173 477
rect 1167 459 1173 465
rect 1167 447 1173 453
rect 1191 471 1197 477
rect 1191 459 1197 465
rect 1191 447 1197 453
rect 1215 471 1221 477
rect 1215 459 1221 465
rect 1215 447 1221 453
rect 1239 471 1245 477
rect 1239 459 1245 465
rect 1239 447 1245 453
rect 1263 471 1269 477
rect 1263 459 1269 465
rect 1263 447 1269 453
rect 1287 471 1293 477
rect 1287 459 1293 465
rect 1287 447 1293 453
rect 1311 471 1317 477
rect 1311 459 1317 465
rect 1311 447 1317 453
rect 1335 471 1341 477
rect 1335 459 1341 465
rect 1335 447 1341 453
rect 1359 471 1365 477
rect 1359 459 1365 465
rect 1359 447 1365 453
rect 1383 471 1389 477
rect 1383 459 1389 465
rect 1383 447 1389 453
rect 1407 471 1413 477
rect 1407 459 1413 465
rect 1407 447 1413 453
rect 1431 471 1437 477
rect 1431 459 1437 465
rect 1431 447 1437 453
rect 1455 471 1461 477
rect 1455 459 1461 465
rect 1455 447 1461 453
rect 1479 471 1485 477
rect 1479 459 1485 465
rect 1479 447 1485 453
<< psubdiff >>
rect -48 213 1524 216
rect -48 207 -45 213
rect -39 207 -33 213
rect -27 207 -21 213
rect -15 207 -9 213
rect -3 207 3 213
rect 9 207 15 213
rect 21 207 27 213
rect 33 207 39 213
rect 45 207 51 213
rect 57 207 63 213
rect 69 207 75 213
rect 81 207 87 213
rect 93 207 99 213
rect 105 207 111 213
rect 117 207 123 213
rect 129 207 135 213
rect 141 207 147 213
rect 153 207 159 213
rect 165 207 171 213
rect 177 207 183 213
rect 189 207 195 213
rect 201 207 207 213
rect 213 207 219 213
rect 225 207 231 213
rect 237 207 243 213
rect 249 207 255 213
rect 261 207 267 213
rect 273 207 279 213
rect 285 207 291 213
rect 297 207 303 213
rect 309 207 315 213
rect 321 207 327 213
rect 333 207 339 213
rect 345 207 351 213
rect 357 207 363 213
rect 369 207 375 213
rect 381 207 387 213
rect 393 207 399 213
rect 405 207 411 213
rect 417 207 423 213
rect 429 207 435 213
rect 441 207 447 213
rect 453 207 459 213
rect 465 207 471 213
rect 477 207 483 213
rect 489 207 495 213
rect 501 207 507 213
rect 513 207 519 213
rect 525 207 531 213
rect 537 207 543 213
rect 549 207 555 213
rect 561 207 567 213
rect 573 207 579 213
rect 585 207 591 213
rect 597 207 603 213
rect 609 207 615 213
rect 621 207 627 213
rect 633 207 639 213
rect 645 207 651 213
rect 657 207 663 213
rect 669 207 675 213
rect 681 207 687 213
rect 693 207 699 213
rect 705 207 711 213
rect 717 207 723 213
rect 729 207 735 213
rect 741 207 747 213
rect 753 207 759 213
rect 765 207 771 213
rect 777 207 783 213
rect 789 207 795 213
rect 801 207 807 213
rect 813 207 819 213
rect 825 207 831 213
rect 837 207 843 213
rect 849 207 855 213
rect 861 207 867 213
rect 873 207 879 213
rect 885 207 891 213
rect 897 207 903 213
rect 909 207 915 213
rect 921 207 927 213
rect 933 207 939 213
rect 945 207 951 213
rect 957 207 963 213
rect 969 207 975 213
rect 981 207 987 213
rect 993 207 999 213
rect 1005 207 1011 213
rect 1017 207 1023 213
rect 1029 207 1035 213
rect 1041 207 1047 213
rect 1053 207 1059 213
rect 1065 207 1071 213
rect 1077 207 1083 213
rect 1089 207 1095 213
rect 1101 207 1107 213
rect 1113 207 1119 213
rect 1125 207 1131 213
rect 1137 207 1143 213
rect 1149 207 1155 213
rect 1161 207 1167 213
rect 1173 207 1179 213
rect 1185 207 1191 213
rect 1197 207 1203 213
rect 1209 207 1215 213
rect 1221 207 1227 213
rect 1233 207 1239 213
rect 1245 207 1251 213
rect 1257 207 1263 213
rect 1269 207 1275 213
rect 1281 207 1287 213
rect 1293 207 1299 213
rect 1305 207 1311 213
rect 1317 207 1323 213
rect 1329 207 1335 213
rect 1341 207 1347 213
rect 1353 207 1359 213
rect 1365 207 1371 213
rect 1377 207 1383 213
rect 1389 207 1395 213
rect 1401 207 1407 213
rect 1413 207 1419 213
rect 1425 207 1431 213
rect 1437 207 1443 213
rect 1449 207 1455 213
rect 1461 207 1467 213
rect 1473 207 1479 213
rect 1485 207 1491 213
rect 1497 207 1503 213
rect 1509 207 1515 213
rect 1521 207 1524 213
rect -48 204 1524 207
rect -48 93 1524 96
rect -48 87 -45 93
rect -39 87 -33 93
rect -27 87 -21 93
rect -15 87 -9 93
rect -3 87 3 93
rect 9 87 15 93
rect 21 87 27 93
rect 33 87 39 93
rect 45 87 51 93
rect 57 87 63 93
rect 69 87 75 93
rect 81 87 87 93
rect 93 87 99 93
rect 105 87 111 93
rect 117 87 123 93
rect 129 87 135 93
rect 141 87 147 93
rect 153 87 159 93
rect 165 87 171 93
rect 177 87 183 93
rect 189 87 195 93
rect 201 87 207 93
rect 213 87 219 93
rect 225 87 231 93
rect 237 87 243 93
rect 249 87 255 93
rect 261 87 267 93
rect 273 87 279 93
rect 285 87 291 93
rect 297 87 303 93
rect 309 87 315 93
rect 321 87 327 93
rect 333 87 339 93
rect 345 87 351 93
rect 357 87 363 93
rect 369 87 375 93
rect 381 87 387 93
rect 393 87 399 93
rect 405 87 411 93
rect 417 87 423 93
rect 429 87 435 93
rect 441 87 447 93
rect 453 87 459 93
rect 465 87 471 93
rect 477 87 483 93
rect 489 87 495 93
rect 501 87 507 93
rect 513 87 519 93
rect 525 87 531 93
rect 537 87 543 93
rect 549 87 555 93
rect 561 87 567 93
rect 573 87 579 93
rect 585 87 591 93
rect 597 87 603 93
rect 609 87 615 93
rect 621 87 627 93
rect 633 87 639 93
rect 645 87 651 93
rect 657 87 663 93
rect 669 87 675 93
rect 681 87 687 93
rect 693 87 699 93
rect 705 87 711 93
rect 717 87 723 93
rect 729 87 735 93
rect 741 87 747 93
rect 753 87 759 93
rect 765 87 771 93
rect 777 87 783 93
rect 789 87 795 93
rect 801 87 807 93
rect 813 87 819 93
rect 825 87 831 93
rect 837 87 843 93
rect 849 87 855 93
rect 861 87 867 93
rect 873 87 879 93
rect 885 87 891 93
rect 897 87 903 93
rect 909 87 915 93
rect 921 87 927 93
rect 933 87 939 93
rect 945 87 951 93
rect 957 87 963 93
rect 969 87 975 93
rect 981 87 987 93
rect 993 87 999 93
rect 1005 87 1011 93
rect 1017 87 1023 93
rect 1029 87 1035 93
rect 1041 87 1047 93
rect 1053 87 1059 93
rect 1065 87 1071 93
rect 1077 87 1083 93
rect 1089 87 1095 93
rect 1101 87 1107 93
rect 1113 87 1119 93
rect 1125 87 1131 93
rect 1137 87 1143 93
rect 1149 87 1155 93
rect 1161 87 1167 93
rect 1173 87 1179 93
rect 1185 87 1191 93
rect 1197 87 1203 93
rect 1209 87 1215 93
rect 1221 87 1227 93
rect 1233 87 1239 93
rect 1245 87 1251 93
rect 1257 87 1263 93
rect 1269 87 1275 93
rect 1281 87 1287 93
rect 1293 87 1299 93
rect 1305 87 1311 93
rect 1317 87 1323 93
rect 1329 87 1335 93
rect 1341 87 1347 93
rect 1353 87 1359 93
rect 1365 87 1371 93
rect 1377 87 1383 93
rect 1389 87 1395 93
rect 1401 87 1407 93
rect 1413 87 1419 93
rect 1425 87 1431 93
rect 1437 87 1443 93
rect 1449 87 1455 93
rect 1461 87 1467 93
rect 1473 87 1479 93
rect 1485 87 1491 93
rect 1497 87 1503 93
rect 1509 87 1515 93
rect 1521 87 1524 93
rect -48 84 1524 87
rect -48 -3 1524 0
rect -48 -9 -45 -3
rect -39 -9 -33 -3
rect -27 -9 -21 -3
rect -15 -9 -9 -3
rect -3 -9 3 -3
rect 9 -9 15 -3
rect 21 -9 27 -3
rect 33 -9 39 -3
rect 45 -9 51 -3
rect 57 -9 63 -3
rect 69 -9 75 -3
rect 81 -9 87 -3
rect 93 -9 99 -3
rect 105 -9 111 -3
rect 117 -9 123 -3
rect 129 -9 135 -3
rect 141 -9 147 -3
rect 153 -9 159 -3
rect 165 -9 171 -3
rect 177 -9 183 -3
rect 189 -9 195 -3
rect 201 -9 207 -3
rect 213 -9 219 -3
rect 225 -9 231 -3
rect 237 -9 243 -3
rect 249 -9 255 -3
rect 261 -9 267 -3
rect 273 -9 279 -3
rect 285 -9 291 -3
rect 297 -9 303 -3
rect 309 -9 315 -3
rect 321 -9 327 -3
rect 333 -9 339 -3
rect 345 -9 351 -3
rect 357 -9 363 -3
rect 369 -9 375 -3
rect 381 -9 387 -3
rect 393 -9 399 -3
rect 405 -9 411 -3
rect 417 -9 423 -3
rect 429 -9 435 -3
rect 441 -9 447 -3
rect 453 -9 459 -3
rect 465 -9 471 -3
rect 477 -9 483 -3
rect 489 -9 495 -3
rect 501 -9 507 -3
rect 513 -9 519 -3
rect 525 -9 531 -3
rect 537 -9 543 -3
rect 549 -9 555 -3
rect 561 -9 567 -3
rect 573 -9 579 -3
rect 585 -9 591 -3
rect 597 -9 603 -3
rect 609 -9 615 -3
rect 621 -9 627 -3
rect 633 -9 639 -3
rect 645 -9 651 -3
rect 657 -9 663 -3
rect 669 -9 675 -3
rect 681 -9 687 -3
rect 693 -9 699 -3
rect 705 -9 711 -3
rect 717 -9 723 -3
rect 729 -9 735 -3
rect 741 -9 747 -3
rect 753 -9 759 -3
rect 765 -9 771 -3
rect 777 -9 783 -3
rect 789 -9 795 -3
rect 801 -9 807 -3
rect 813 -9 819 -3
rect 825 -9 831 -3
rect 837 -9 843 -3
rect 849 -9 855 -3
rect 861 -9 867 -3
rect 873 -9 879 -3
rect 885 -9 891 -3
rect 897 -9 903 -3
rect 909 -9 915 -3
rect 921 -9 927 -3
rect 933 -9 939 -3
rect 945 -9 951 -3
rect 957 -9 963 -3
rect 969 -9 975 -3
rect 981 -9 987 -3
rect 993 -9 999 -3
rect 1005 -9 1011 -3
rect 1017 -9 1023 -3
rect 1029 -9 1035 -3
rect 1041 -9 1047 -3
rect 1053 -9 1059 -3
rect 1065 -9 1071 -3
rect 1077 -9 1083 -3
rect 1089 -9 1095 -3
rect 1101 -9 1107 -3
rect 1113 -9 1119 -3
rect 1125 -9 1131 -3
rect 1137 -9 1143 -3
rect 1149 -9 1155 -3
rect 1161 -9 1167 -3
rect 1173 -9 1179 -3
rect 1185 -9 1191 -3
rect 1197 -9 1203 -3
rect 1209 -9 1215 -3
rect 1221 -9 1227 -3
rect 1233 -9 1239 -3
rect 1245 -9 1251 -3
rect 1257 -9 1263 -3
rect 1269 -9 1275 -3
rect 1281 -9 1287 -3
rect 1293 -9 1299 -3
rect 1305 -9 1311 -3
rect 1317 -9 1323 -3
rect 1329 -9 1335 -3
rect 1341 -9 1347 -3
rect 1353 -9 1359 -3
rect 1365 -9 1371 -3
rect 1377 -9 1383 -3
rect 1389 -9 1395 -3
rect 1401 -9 1407 -3
rect 1413 -9 1419 -3
rect 1425 -9 1431 -3
rect 1437 -9 1443 -3
rect 1449 -9 1455 -3
rect 1461 -9 1467 -3
rect 1473 -9 1479 -3
rect 1485 -9 1491 -3
rect 1497 -9 1503 -3
rect 1509 -9 1515 -3
rect 1521 -9 1524 -3
rect -48 -12 1524 -9
<< mvpsubdiff >>
rect -60 621 1536 624
rect -60 615 -57 621
rect -51 615 -45 621
rect -39 615 -33 621
rect -27 615 -21 621
rect -15 615 -9 621
rect -3 615 3 621
rect 9 615 15 621
rect 21 615 27 621
rect 33 615 39 621
rect 45 615 51 621
rect 57 615 63 621
rect 69 615 75 621
rect 81 615 87 621
rect 93 615 99 621
rect 105 615 111 621
rect 117 615 123 621
rect 129 615 135 621
rect 141 615 147 621
rect 153 615 159 621
rect 165 615 171 621
rect 177 615 183 621
rect 189 615 195 621
rect 201 615 207 621
rect 213 615 219 621
rect 225 615 231 621
rect 237 615 243 621
rect 249 615 255 621
rect 261 615 267 621
rect 273 615 279 621
rect 285 615 291 621
rect 297 615 303 621
rect 309 615 315 621
rect 321 615 327 621
rect 333 615 339 621
rect 345 615 351 621
rect 357 615 363 621
rect 369 615 375 621
rect 381 615 387 621
rect 393 615 399 621
rect 405 615 411 621
rect 417 615 423 621
rect 429 615 435 621
rect 441 615 447 621
rect 453 615 459 621
rect 465 615 471 621
rect 477 615 483 621
rect 489 615 495 621
rect 501 615 507 621
rect 513 615 519 621
rect 525 615 531 621
rect 537 615 543 621
rect 549 615 555 621
rect 561 615 567 621
rect 573 615 579 621
rect 585 615 591 621
rect 597 615 603 621
rect 609 615 615 621
rect 621 615 627 621
rect 633 615 639 621
rect 645 615 651 621
rect 657 615 663 621
rect 669 615 675 621
rect 681 615 687 621
rect 693 615 699 621
rect 705 615 711 621
rect 717 615 723 621
rect 729 615 735 621
rect 741 615 747 621
rect 753 615 759 621
rect 765 615 771 621
rect 777 615 783 621
rect 789 615 795 621
rect 801 615 807 621
rect 813 615 819 621
rect 825 615 831 621
rect 837 615 843 621
rect 849 615 855 621
rect 861 615 867 621
rect 873 615 879 621
rect 885 615 891 621
rect 897 615 903 621
rect 909 615 915 621
rect 921 615 927 621
rect 933 615 939 621
rect 945 615 951 621
rect 957 615 963 621
rect 969 615 975 621
rect 981 615 987 621
rect 993 615 999 621
rect 1005 615 1011 621
rect 1017 615 1023 621
rect 1029 615 1035 621
rect 1041 615 1047 621
rect 1053 615 1059 621
rect 1065 615 1071 621
rect 1077 615 1083 621
rect 1089 615 1095 621
rect 1101 615 1107 621
rect 1113 615 1119 621
rect 1125 615 1131 621
rect 1137 615 1143 621
rect 1149 615 1155 621
rect 1161 615 1167 621
rect 1173 615 1179 621
rect 1185 615 1191 621
rect 1197 615 1203 621
rect 1209 615 1215 621
rect 1221 615 1227 621
rect 1233 615 1239 621
rect 1245 615 1251 621
rect 1257 615 1263 621
rect 1269 615 1275 621
rect 1281 615 1287 621
rect 1293 615 1299 621
rect 1305 615 1311 621
rect 1317 615 1323 621
rect 1329 615 1335 621
rect 1341 615 1347 621
rect 1353 615 1359 621
rect 1365 615 1371 621
rect 1377 615 1383 621
rect 1389 615 1395 621
rect 1401 615 1407 621
rect 1413 615 1419 621
rect 1425 615 1431 621
rect 1437 615 1443 621
rect 1449 615 1455 621
rect 1461 615 1467 621
rect 1473 615 1479 621
rect 1485 615 1491 621
rect 1497 615 1503 621
rect 1509 615 1515 621
rect 1521 615 1527 621
rect 1533 615 1536 621
rect -60 612 1536 615
rect -60 609 -48 612
rect -60 603 -57 609
rect -51 603 -48 609
rect -60 597 -48 603
rect 1524 609 1536 612
rect 1524 603 1527 609
rect 1533 603 1536 609
rect -60 591 -57 597
rect -51 591 -48 597
rect -60 585 -48 591
rect -60 579 -57 585
rect -51 579 -48 585
rect -60 573 -48 579
rect -60 567 -57 573
rect -51 567 -48 573
rect -60 561 -48 567
rect -60 555 -57 561
rect -51 555 -48 561
rect -60 549 -48 555
rect -60 543 -57 549
rect -51 543 -48 549
rect -60 537 -48 543
rect -60 531 -57 537
rect -51 531 -48 537
rect -60 525 -48 531
rect -60 519 -57 525
rect -51 519 -48 525
rect -60 513 -48 519
rect -60 507 -57 513
rect -51 507 -48 513
rect -60 501 -48 507
rect -60 495 -57 501
rect -51 495 -48 501
rect -60 489 -48 495
rect -60 483 -57 489
rect -51 483 -48 489
rect -60 477 -48 483
rect -60 471 -57 477
rect -51 471 -48 477
rect -60 465 -48 471
rect -60 459 -57 465
rect -51 459 -48 465
rect -60 453 -48 459
rect -60 447 -57 453
rect -51 447 -48 453
rect -60 441 -48 447
rect -60 435 -57 441
rect -51 435 -48 441
rect -60 429 -48 435
rect -60 423 -57 429
rect -51 423 -48 429
rect -60 417 -48 423
rect -60 411 -57 417
rect -51 411 -48 417
rect -60 405 -48 411
rect -60 399 -57 405
rect -51 399 -48 405
rect -60 393 -48 399
rect -60 387 -57 393
rect -51 387 -48 393
rect -60 381 -48 387
rect -60 375 -57 381
rect -51 375 -48 381
rect -60 369 -48 375
rect -60 363 -57 369
rect -51 363 -48 369
rect -60 357 -48 363
rect -60 351 -57 357
rect -51 351 -48 357
rect -60 345 -48 351
rect 1524 597 1536 603
rect 1524 591 1527 597
rect 1533 591 1536 597
rect 1524 585 1536 591
rect 1524 579 1527 585
rect 1533 579 1536 585
rect 1524 573 1536 579
rect 1524 567 1527 573
rect 1533 567 1536 573
rect 1524 561 1536 567
rect 1524 555 1527 561
rect 1533 555 1536 561
rect 1524 549 1536 555
rect 1524 543 1527 549
rect 1533 543 1536 549
rect 1524 537 1536 543
rect 1524 531 1527 537
rect 1533 531 1536 537
rect 1524 525 1536 531
rect 1524 519 1527 525
rect 1533 519 1536 525
rect 1524 513 1536 519
rect 1524 507 1527 513
rect 1533 507 1536 513
rect 1524 501 1536 507
rect 1524 495 1527 501
rect 1533 495 1536 501
rect 1524 489 1536 495
rect 1524 483 1527 489
rect 1533 483 1536 489
rect 1524 477 1536 483
rect 1524 471 1527 477
rect 1533 471 1536 477
rect 1524 465 1536 471
rect 1524 459 1527 465
rect 1533 459 1536 465
rect 1524 453 1536 459
rect 1524 447 1527 453
rect 1533 447 1536 453
rect 1524 441 1536 447
rect 1524 435 1527 441
rect 1533 435 1536 441
rect 1524 429 1536 435
rect 1524 423 1527 429
rect 1533 423 1536 429
rect 1524 417 1536 423
rect 1524 411 1527 417
rect 1533 411 1536 417
rect 1524 405 1536 411
rect 1524 399 1527 405
rect 1533 399 1536 405
rect 1524 393 1536 399
rect 1524 387 1527 393
rect 1533 387 1536 393
rect 1524 381 1536 387
rect 1524 375 1527 381
rect 1533 375 1536 381
rect 1524 369 1536 375
rect 1524 363 1527 369
rect 1533 363 1536 369
rect 1524 357 1536 363
rect 1524 351 1527 357
rect 1533 351 1536 357
rect -60 339 -57 345
rect -51 339 -48 345
rect -60 336 -48 339
rect 1524 345 1536 351
rect 1524 339 1527 345
rect 1533 339 1536 345
rect 1524 336 1536 339
rect -60 333 1536 336
rect -60 327 -57 333
rect -51 327 -45 333
rect -39 327 -33 333
rect -27 327 -21 333
rect -15 327 -9 333
rect -3 327 3 333
rect 9 327 15 333
rect 21 327 27 333
rect 33 327 39 333
rect 45 327 51 333
rect 57 327 63 333
rect 69 327 75 333
rect 81 327 87 333
rect 93 327 99 333
rect 105 327 111 333
rect 117 327 123 333
rect 129 327 135 333
rect 141 327 147 333
rect 153 327 159 333
rect 165 327 171 333
rect 177 327 183 333
rect 189 327 195 333
rect 201 327 207 333
rect 213 327 219 333
rect 225 327 231 333
rect 237 327 243 333
rect 249 327 255 333
rect 261 327 267 333
rect 273 327 279 333
rect 285 327 291 333
rect 297 327 303 333
rect 309 327 315 333
rect 321 327 327 333
rect 333 327 339 333
rect 345 327 351 333
rect 357 327 363 333
rect 369 327 375 333
rect 381 327 387 333
rect 393 327 399 333
rect 405 327 411 333
rect 417 327 423 333
rect 429 327 435 333
rect 441 327 447 333
rect 453 327 459 333
rect 465 327 471 333
rect 477 327 483 333
rect 489 327 495 333
rect 501 327 507 333
rect 513 327 519 333
rect 525 327 531 333
rect 537 327 543 333
rect 549 327 555 333
rect 561 327 567 333
rect 573 327 579 333
rect 585 327 591 333
rect 597 327 603 333
rect 609 327 615 333
rect 621 327 627 333
rect 633 327 639 333
rect 645 327 651 333
rect 657 327 663 333
rect 669 327 675 333
rect 681 327 687 333
rect 693 327 699 333
rect 705 327 711 333
rect 717 327 723 333
rect 729 327 735 333
rect 741 327 747 333
rect 753 327 759 333
rect 765 327 771 333
rect 777 327 783 333
rect 789 327 795 333
rect 801 327 807 333
rect 813 327 819 333
rect 825 327 831 333
rect 837 327 843 333
rect 849 327 855 333
rect 861 327 867 333
rect 873 327 879 333
rect 885 327 891 333
rect 897 327 903 333
rect 909 327 915 333
rect 921 327 927 333
rect 933 327 939 333
rect 945 327 951 333
rect 957 327 963 333
rect 969 327 975 333
rect 981 327 987 333
rect 993 327 999 333
rect 1005 327 1011 333
rect 1017 327 1023 333
rect 1029 327 1035 333
rect 1041 327 1047 333
rect 1053 327 1059 333
rect 1065 327 1071 333
rect 1077 327 1083 333
rect 1089 327 1095 333
rect 1101 327 1107 333
rect 1113 327 1119 333
rect 1125 327 1131 333
rect 1137 327 1143 333
rect 1149 327 1155 333
rect 1161 327 1167 333
rect 1173 327 1179 333
rect 1185 327 1191 333
rect 1197 327 1203 333
rect 1209 327 1215 333
rect 1221 327 1227 333
rect 1233 327 1239 333
rect 1245 327 1251 333
rect 1257 327 1263 333
rect 1269 327 1275 333
rect 1281 327 1287 333
rect 1293 327 1299 333
rect 1305 327 1311 333
rect 1317 327 1323 333
rect 1329 327 1335 333
rect 1341 327 1347 333
rect 1353 327 1359 333
rect 1365 327 1371 333
rect 1377 327 1383 333
rect 1389 327 1395 333
rect 1401 327 1407 333
rect 1413 327 1419 333
rect 1425 327 1431 333
rect 1437 327 1443 333
rect 1449 327 1455 333
rect 1461 327 1467 333
rect 1473 327 1479 333
rect 1485 327 1491 333
rect 1497 327 1503 333
rect 1509 327 1515 333
rect 1521 327 1527 333
rect 1533 327 1536 333
rect -60 324 1536 327
rect -60 321 -48 324
rect -60 315 -57 321
rect -51 315 -48 321
rect -60 309 -48 315
rect 1524 321 1536 324
rect 1524 315 1527 321
rect 1533 315 1536 321
rect -60 303 -57 309
rect -51 303 -48 309
rect -60 297 -48 303
rect -60 291 -57 297
rect -51 291 -48 297
rect -60 285 -48 291
rect 1524 309 1536 315
rect 1524 303 1527 309
rect 1533 303 1536 309
rect 1524 297 1536 303
rect 1524 291 1527 297
rect 1533 291 1536 297
rect -60 279 -57 285
rect -51 279 -48 285
rect -60 273 -48 279
rect -60 267 -57 273
rect -51 267 -48 273
rect -60 261 -48 267
rect -60 255 -57 261
rect -51 255 -48 261
rect -60 249 -48 255
rect 1524 285 1536 291
rect 1524 279 1527 285
rect 1533 279 1536 285
rect 1524 273 1536 279
rect 1524 267 1527 273
rect 1533 267 1536 273
rect 1524 261 1536 267
rect 1524 255 1527 261
rect 1533 255 1536 261
rect -60 243 -57 249
rect -51 243 -48 249
rect 1524 249 1536 255
rect -60 237 -48 243
rect -60 231 -57 237
rect -51 231 -48 237
rect -60 225 -48 231
rect -60 219 -57 225
rect -51 219 -48 225
rect -60 213 -48 219
rect 1524 243 1527 249
rect 1533 243 1536 249
rect 1524 237 1536 243
rect 1524 231 1527 237
rect 1533 231 1536 237
rect 1524 225 1536 231
rect 1524 219 1527 225
rect 1533 219 1536 225
rect 1524 213 1536 219
rect -60 207 -57 213
rect -51 207 -48 213
rect 1524 207 1527 213
rect 1533 207 1536 213
rect -60 201 -48 207
rect -60 195 -57 201
rect -51 195 -48 201
rect -60 189 -48 195
rect -60 183 -57 189
rect -51 183 -48 189
rect -60 177 -48 183
rect -60 171 -57 177
rect -51 171 -48 177
rect -60 165 -48 171
rect -60 159 -57 165
rect -51 159 -48 165
rect -60 153 -48 159
rect -60 147 -57 153
rect -51 147 -48 153
rect -60 141 -48 147
rect -60 135 -57 141
rect -51 135 -48 141
rect -60 129 -48 135
rect -60 123 -57 129
rect -51 123 -48 129
rect -60 117 -48 123
rect -60 111 -57 117
rect -51 111 -48 117
rect -60 105 -48 111
rect -60 99 -57 105
rect -51 99 -48 105
rect -60 93 -48 99
rect 1524 201 1536 207
rect 1524 195 1527 201
rect 1533 195 1536 201
rect 1524 189 1536 195
rect 1524 183 1527 189
rect 1533 183 1536 189
rect 1524 177 1536 183
rect 1524 171 1527 177
rect 1533 171 1536 177
rect 1524 165 1536 171
rect 1524 159 1527 165
rect 1533 159 1536 165
rect 1524 153 1536 159
rect 1524 147 1527 153
rect 1533 147 1536 153
rect 1524 141 1536 147
rect 1524 135 1527 141
rect 1533 135 1536 141
rect 1524 129 1536 135
rect 1524 123 1527 129
rect 1533 123 1536 129
rect 1524 117 1536 123
rect 1524 111 1527 117
rect 1533 111 1536 117
rect 1524 105 1536 111
rect 1524 99 1527 105
rect 1533 99 1536 105
rect 1524 93 1536 99
rect -60 87 -57 93
rect -51 87 -48 93
rect 1524 87 1527 93
rect 1533 87 1536 93
rect -60 81 -48 87
rect -60 75 -57 81
rect -51 75 -48 81
rect -60 69 -48 75
rect 1524 81 1536 87
rect 1524 75 1527 81
rect 1533 75 1536 81
rect -60 63 -57 69
rect -51 63 -48 69
rect -60 57 -48 63
rect -60 51 -57 57
rect -51 51 -48 57
rect -60 45 -48 51
rect 1524 69 1536 75
rect 1524 63 1527 69
rect 1533 63 1536 69
rect 1524 57 1536 63
rect 1524 51 1527 57
rect 1533 51 1536 57
rect -60 39 -57 45
rect -51 39 -48 45
rect -60 33 -48 39
rect -60 27 -57 33
rect -51 27 -48 33
rect -60 21 -48 27
rect -60 15 -57 21
rect -51 15 -48 21
rect -60 9 -48 15
rect 1524 45 1536 51
rect 1524 39 1527 45
rect 1533 39 1536 45
rect 1524 33 1536 39
rect 1524 27 1527 33
rect 1533 27 1536 33
rect 1524 21 1536 27
rect 1524 15 1527 21
rect 1533 15 1536 21
rect -60 3 -57 9
rect -51 3 -48 9
rect 1524 9 1536 15
rect -60 -3 -48 3
rect 1524 3 1527 9
rect 1533 3 1536 9
rect 1524 -3 1536 3
rect -60 -9 -57 -3
rect -51 -9 -48 -3
rect 1524 -9 1527 -3
rect 1533 -9 1536 -3
rect -60 -12 -48 -9
rect 1524 -12 1536 -9
<< mvnsubdiff >>
rect -36 597 1512 600
rect -36 591 -33 597
rect -27 591 -21 597
rect -15 591 -9 597
rect -3 591 3 597
rect 9 591 15 597
rect 21 591 27 597
rect 33 591 39 597
rect 45 591 51 597
rect 57 591 63 597
rect 69 591 75 597
rect 81 591 87 597
rect 93 591 99 597
rect 105 591 111 597
rect 117 591 123 597
rect 129 591 135 597
rect 141 591 147 597
rect 153 591 159 597
rect 165 591 171 597
rect 177 591 183 597
rect 189 591 195 597
rect 201 591 207 597
rect 213 591 219 597
rect 225 591 231 597
rect 237 591 243 597
rect 249 591 255 597
rect 261 591 267 597
rect 273 591 279 597
rect 285 591 291 597
rect 297 591 303 597
rect 309 591 315 597
rect 321 591 327 597
rect 333 591 339 597
rect 345 591 351 597
rect 357 591 363 597
rect 369 591 375 597
rect 381 591 387 597
rect 393 591 399 597
rect 405 591 411 597
rect 417 591 423 597
rect 429 591 435 597
rect 441 591 447 597
rect 453 591 459 597
rect 465 591 471 597
rect 477 591 483 597
rect 489 591 495 597
rect 501 591 507 597
rect 513 591 519 597
rect 525 591 531 597
rect 537 591 543 597
rect 549 591 555 597
rect 561 591 567 597
rect 573 591 579 597
rect 585 591 591 597
rect 597 591 603 597
rect 609 591 615 597
rect 621 591 627 597
rect 633 591 639 597
rect 645 591 651 597
rect 657 591 663 597
rect 669 591 675 597
rect 681 591 687 597
rect 693 591 699 597
rect 705 591 711 597
rect 717 591 723 597
rect 729 591 735 597
rect 741 591 747 597
rect 753 591 759 597
rect 765 591 771 597
rect 777 591 783 597
rect 789 591 795 597
rect 801 591 807 597
rect 813 591 819 597
rect 825 591 831 597
rect 837 591 843 597
rect 849 591 855 597
rect 861 591 867 597
rect 873 591 879 597
rect 885 591 891 597
rect 897 591 903 597
rect 909 591 915 597
rect 921 591 927 597
rect 933 591 939 597
rect 945 591 951 597
rect 957 591 963 597
rect 969 591 975 597
rect 981 591 987 597
rect 993 591 999 597
rect 1005 591 1011 597
rect 1017 591 1023 597
rect 1029 591 1035 597
rect 1041 591 1047 597
rect 1053 591 1059 597
rect 1065 591 1071 597
rect 1077 591 1083 597
rect 1089 591 1095 597
rect 1101 591 1107 597
rect 1113 591 1119 597
rect 1125 591 1131 597
rect 1137 591 1143 597
rect 1149 591 1155 597
rect 1161 591 1167 597
rect 1173 591 1179 597
rect 1185 591 1191 597
rect 1197 591 1203 597
rect 1209 591 1215 597
rect 1221 591 1227 597
rect 1233 591 1239 597
rect 1245 591 1251 597
rect 1257 591 1263 597
rect 1269 591 1275 597
rect 1281 591 1287 597
rect 1293 591 1299 597
rect 1305 591 1311 597
rect 1317 591 1323 597
rect 1329 591 1335 597
rect 1341 591 1347 597
rect 1353 591 1359 597
rect 1365 591 1371 597
rect 1377 591 1383 597
rect 1389 591 1395 597
rect 1401 591 1407 597
rect 1413 591 1419 597
rect 1425 591 1431 597
rect 1437 591 1443 597
rect 1449 591 1455 597
rect 1461 591 1467 597
rect 1473 591 1479 597
rect 1485 591 1491 597
rect 1497 591 1503 597
rect 1509 591 1512 597
rect -36 588 1512 591
rect -36 585 -24 588
rect -36 579 -33 585
rect -27 579 -24 585
rect 1500 585 1512 588
rect -36 573 -24 579
rect 1500 579 1503 585
rect 1509 579 1512 585
rect -36 567 -33 573
rect -27 567 -24 573
rect -36 561 -24 567
rect -36 555 -33 561
rect -27 555 -24 561
rect -36 549 -24 555
rect -36 543 -33 549
rect -27 543 -24 549
rect -36 537 -24 543
rect 1500 573 1512 579
rect 1500 567 1503 573
rect 1509 567 1512 573
rect 1500 561 1512 567
rect 1500 555 1503 561
rect 1509 555 1512 561
rect 1500 549 1512 555
rect 1500 543 1503 549
rect 1509 543 1512 549
rect -36 531 -33 537
rect -27 531 -24 537
rect -36 525 -24 531
rect -36 519 -33 525
rect -27 519 -24 525
rect -36 513 -24 519
rect 1500 537 1512 543
rect 1500 531 1503 537
rect 1509 531 1512 537
rect 1500 525 1512 531
rect 1500 519 1503 525
rect 1509 519 1512 525
rect -36 507 -33 513
rect -27 507 -24 513
rect -36 504 -24 507
rect 1500 513 1512 519
rect 1500 507 1503 513
rect 1509 507 1512 513
rect 1500 504 1512 507
rect -36 501 1512 504
rect -36 495 -33 501
rect -27 495 -21 501
rect -15 495 -9 501
rect -3 495 3 501
rect 9 495 15 501
rect 21 495 27 501
rect 33 495 39 501
rect 45 495 51 501
rect 57 495 63 501
rect 69 495 75 501
rect 81 495 87 501
rect 93 495 99 501
rect 105 495 111 501
rect 117 495 123 501
rect 129 495 135 501
rect 141 495 147 501
rect 153 495 159 501
rect 165 495 171 501
rect 177 495 183 501
rect 189 495 195 501
rect 201 495 207 501
rect 213 495 219 501
rect 225 495 231 501
rect 237 495 243 501
rect 249 495 255 501
rect 261 495 267 501
rect 273 495 279 501
rect 285 495 291 501
rect 297 495 303 501
rect 309 495 315 501
rect 321 495 327 501
rect 333 495 339 501
rect 345 495 351 501
rect 357 495 363 501
rect 369 495 375 501
rect 381 495 387 501
rect 393 495 399 501
rect 405 495 411 501
rect 417 495 423 501
rect 429 495 435 501
rect 441 495 447 501
rect 453 495 459 501
rect 465 495 471 501
rect 477 495 483 501
rect 489 495 495 501
rect 501 495 507 501
rect 513 495 519 501
rect 525 495 531 501
rect 537 495 543 501
rect 549 495 555 501
rect 561 495 567 501
rect 573 495 579 501
rect 585 495 591 501
rect 597 495 603 501
rect 609 495 615 501
rect 621 495 627 501
rect 633 495 639 501
rect 645 495 651 501
rect 657 495 663 501
rect 669 495 675 501
rect 681 495 687 501
rect 693 495 699 501
rect 705 495 711 501
rect 717 495 723 501
rect 729 495 735 501
rect 741 495 747 501
rect 753 495 759 501
rect 765 495 771 501
rect 777 495 783 501
rect 789 495 795 501
rect 801 495 807 501
rect 813 495 819 501
rect 825 495 831 501
rect 837 495 843 501
rect 849 495 855 501
rect 861 495 867 501
rect 873 495 879 501
rect 885 495 891 501
rect 897 495 903 501
rect 909 495 915 501
rect 921 495 927 501
rect 933 495 939 501
rect 945 495 951 501
rect 957 495 963 501
rect 969 495 975 501
rect 981 495 987 501
rect 993 495 999 501
rect 1005 495 1011 501
rect 1017 495 1023 501
rect 1029 495 1035 501
rect 1041 495 1047 501
rect 1053 495 1059 501
rect 1065 495 1071 501
rect 1077 495 1083 501
rect 1089 495 1095 501
rect 1101 495 1107 501
rect 1113 495 1119 501
rect 1125 495 1131 501
rect 1137 495 1143 501
rect 1149 495 1155 501
rect 1161 495 1167 501
rect 1173 495 1179 501
rect 1185 495 1191 501
rect 1197 495 1203 501
rect 1209 495 1215 501
rect 1221 495 1227 501
rect 1233 495 1239 501
rect 1245 495 1251 501
rect 1257 495 1263 501
rect 1269 495 1275 501
rect 1281 495 1287 501
rect 1293 495 1299 501
rect 1305 495 1311 501
rect 1317 495 1323 501
rect 1329 495 1335 501
rect 1341 495 1347 501
rect 1353 495 1359 501
rect 1365 495 1371 501
rect 1377 495 1383 501
rect 1389 495 1395 501
rect 1401 495 1407 501
rect 1413 495 1419 501
rect 1425 495 1431 501
rect 1437 495 1443 501
rect 1449 495 1455 501
rect 1461 495 1467 501
rect 1473 495 1479 501
rect 1485 495 1491 501
rect 1497 495 1503 501
rect 1509 495 1512 501
rect -36 492 1512 495
rect -36 489 -24 492
rect -36 483 -33 489
rect -27 483 -24 489
rect 1500 489 1512 492
rect -36 477 -24 483
rect 1500 483 1503 489
rect 1509 483 1512 489
rect -36 471 -33 477
rect -27 471 -24 477
rect -36 465 -24 471
rect -36 459 -33 465
rect -27 459 -24 465
rect -36 453 -24 459
rect -36 447 -33 453
rect -27 447 -24 453
rect -36 441 -24 447
rect 1500 477 1512 483
rect 1500 471 1503 477
rect 1509 471 1512 477
rect 1500 465 1512 471
rect 1500 459 1503 465
rect 1509 459 1512 465
rect 1500 453 1512 459
rect 1500 447 1503 453
rect 1509 447 1512 453
rect -36 435 -33 441
rect -27 435 -24 441
rect -36 429 -24 435
rect -36 423 -33 429
rect -27 423 -24 429
rect -36 417 -24 423
rect 1500 441 1512 447
rect 1500 435 1503 441
rect 1509 435 1512 441
rect 1500 429 1512 435
rect 1500 423 1503 429
rect 1509 423 1512 429
rect -36 411 -33 417
rect -27 411 -24 417
rect -36 408 -24 411
rect 1500 417 1512 423
rect 1500 411 1503 417
rect 1509 411 1512 417
rect 1500 408 1512 411
rect -36 405 1512 408
rect -36 399 -33 405
rect -27 399 -21 405
rect -15 399 -9 405
rect -3 399 3 405
rect 9 399 15 405
rect 21 399 27 405
rect 33 399 39 405
rect 45 399 51 405
rect 57 399 63 405
rect 69 399 75 405
rect 81 399 87 405
rect 93 399 99 405
rect 105 399 111 405
rect 117 399 123 405
rect 129 399 135 405
rect 141 399 147 405
rect 153 399 159 405
rect 165 399 171 405
rect 177 399 183 405
rect 189 399 195 405
rect 201 399 207 405
rect 213 399 219 405
rect 225 399 231 405
rect 237 399 243 405
rect 249 399 255 405
rect 261 399 267 405
rect 273 399 279 405
rect 285 399 291 405
rect 297 399 303 405
rect 309 399 315 405
rect 321 399 327 405
rect 333 399 339 405
rect 345 399 351 405
rect 357 399 363 405
rect 369 399 375 405
rect 381 399 387 405
rect 393 399 399 405
rect 405 399 411 405
rect 417 399 423 405
rect 429 399 435 405
rect 441 399 447 405
rect 453 399 459 405
rect 465 399 471 405
rect 477 399 483 405
rect 489 399 495 405
rect 501 399 507 405
rect 513 399 519 405
rect 525 399 531 405
rect 537 399 543 405
rect 549 399 555 405
rect 561 399 567 405
rect 573 399 579 405
rect 585 399 591 405
rect 597 399 603 405
rect 609 399 615 405
rect 621 399 627 405
rect 633 399 639 405
rect 645 399 651 405
rect 657 399 663 405
rect 669 399 675 405
rect 681 399 687 405
rect 693 399 699 405
rect 705 399 711 405
rect 717 399 723 405
rect 729 399 735 405
rect 741 399 747 405
rect 753 399 759 405
rect 765 399 771 405
rect 777 399 783 405
rect 789 399 795 405
rect 801 399 807 405
rect 813 399 819 405
rect 825 399 831 405
rect 837 399 843 405
rect 849 399 855 405
rect 861 399 867 405
rect 873 399 879 405
rect 885 399 891 405
rect 897 399 903 405
rect 909 399 915 405
rect 921 399 927 405
rect 933 399 939 405
rect 945 399 951 405
rect 957 399 963 405
rect 969 399 975 405
rect 981 399 987 405
rect 993 399 999 405
rect 1005 399 1011 405
rect 1017 399 1023 405
rect 1029 399 1035 405
rect 1041 399 1047 405
rect 1053 399 1059 405
rect 1065 399 1071 405
rect 1077 399 1083 405
rect 1089 399 1095 405
rect 1101 399 1107 405
rect 1113 399 1119 405
rect 1125 399 1131 405
rect 1137 399 1143 405
rect 1149 399 1155 405
rect 1161 399 1167 405
rect 1173 399 1179 405
rect 1185 399 1191 405
rect 1197 399 1203 405
rect 1209 399 1215 405
rect 1221 399 1227 405
rect 1233 399 1239 405
rect 1245 399 1251 405
rect 1257 399 1263 405
rect 1269 399 1275 405
rect 1281 399 1287 405
rect 1293 399 1299 405
rect 1305 399 1311 405
rect 1317 399 1323 405
rect 1329 399 1335 405
rect 1341 399 1347 405
rect 1353 399 1359 405
rect 1365 399 1371 405
rect 1377 399 1383 405
rect 1389 399 1395 405
rect 1401 399 1407 405
rect 1413 399 1419 405
rect 1425 399 1431 405
rect 1437 399 1443 405
rect 1449 399 1455 405
rect 1461 399 1467 405
rect 1473 399 1479 405
rect 1485 399 1491 405
rect 1497 399 1503 405
rect 1509 399 1512 405
rect -36 396 1512 399
rect -36 393 -24 396
rect -36 387 -33 393
rect -27 387 -24 393
rect -36 381 -24 387
rect -36 375 -33 381
rect -27 375 -24 381
rect -36 369 -24 375
rect -36 363 -33 369
rect -27 363 -24 369
rect -36 360 -24 363
rect 1500 393 1512 396
rect 1500 387 1503 393
rect 1509 387 1512 393
rect 1500 381 1512 387
rect 1500 375 1503 381
rect 1509 375 1512 381
rect 1500 369 1512 375
rect 1500 363 1503 369
rect 1509 363 1512 369
rect 1500 360 1512 363
rect -36 357 1512 360
rect -36 351 -33 357
rect -27 351 -21 357
rect -15 351 -9 357
rect -3 351 3 357
rect 9 351 15 357
rect 21 351 27 357
rect 33 351 39 357
rect 45 351 51 357
rect 57 351 63 357
rect 69 351 75 357
rect 81 351 87 357
rect 93 351 99 357
rect 105 351 111 357
rect 117 351 123 357
rect 129 351 135 357
rect 141 351 147 357
rect 153 351 159 357
rect 165 351 171 357
rect 177 351 183 357
rect 189 351 195 357
rect 201 351 207 357
rect 213 351 219 357
rect 225 351 231 357
rect 237 351 243 357
rect 249 351 255 357
rect 261 351 267 357
rect 273 351 279 357
rect 285 351 291 357
rect 297 351 303 357
rect 309 351 315 357
rect 321 351 327 357
rect 333 351 339 357
rect 345 351 351 357
rect 357 351 363 357
rect 369 351 375 357
rect 381 351 387 357
rect 393 351 399 357
rect 405 351 411 357
rect 417 351 423 357
rect 429 351 435 357
rect 441 351 447 357
rect 453 351 459 357
rect 465 351 471 357
rect 477 351 483 357
rect 489 351 495 357
rect 501 351 507 357
rect 513 351 519 357
rect 525 351 531 357
rect 537 351 543 357
rect 549 351 555 357
rect 561 351 567 357
rect 573 351 579 357
rect 585 351 591 357
rect 597 351 603 357
rect 609 351 615 357
rect 621 351 627 357
rect 633 351 639 357
rect 645 351 651 357
rect 657 351 663 357
rect 669 351 675 357
rect 681 351 687 357
rect 693 351 699 357
rect 705 351 711 357
rect 717 351 723 357
rect 729 351 735 357
rect 741 351 747 357
rect 753 351 759 357
rect 765 351 771 357
rect 777 351 783 357
rect 789 351 795 357
rect 801 351 807 357
rect 813 351 819 357
rect 825 351 831 357
rect 837 351 843 357
rect 849 351 855 357
rect 861 351 867 357
rect 873 351 879 357
rect 885 351 891 357
rect 897 351 903 357
rect 909 351 915 357
rect 921 351 927 357
rect 933 351 939 357
rect 945 351 951 357
rect 957 351 963 357
rect 969 351 975 357
rect 981 351 987 357
rect 993 351 999 357
rect 1005 351 1011 357
rect 1017 351 1023 357
rect 1029 351 1035 357
rect 1041 351 1047 357
rect 1053 351 1059 357
rect 1065 351 1071 357
rect 1077 351 1083 357
rect 1089 351 1095 357
rect 1101 351 1107 357
rect 1113 351 1119 357
rect 1125 351 1131 357
rect 1137 351 1143 357
rect 1149 351 1155 357
rect 1161 351 1167 357
rect 1173 351 1179 357
rect 1185 351 1191 357
rect 1197 351 1203 357
rect 1209 351 1215 357
rect 1221 351 1227 357
rect 1233 351 1239 357
rect 1245 351 1251 357
rect 1257 351 1263 357
rect 1269 351 1275 357
rect 1281 351 1287 357
rect 1293 351 1299 357
rect 1305 351 1311 357
rect 1317 351 1323 357
rect 1329 351 1335 357
rect 1341 351 1347 357
rect 1353 351 1359 357
rect 1365 351 1371 357
rect 1377 351 1383 357
rect 1389 351 1395 357
rect 1401 351 1407 357
rect 1413 351 1419 357
rect 1425 351 1431 357
rect 1437 351 1443 357
rect 1449 351 1455 357
rect 1461 351 1467 357
rect 1473 351 1479 357
rect 1485 351 1491 357
rect 1497 351 1503 357
rect 1509 351 1512 357
rect -36 348 1512 351
<< psubdiffcont >>
rect -45 207 -39 213
rect -33 207 -27 213
rect -21 207 -15 213
rect -9 207 -3 213
rect 3 207 9 213
rect 15 207 21 213
rect 27 207 33 213
rect 39 207 45 213
rect 51 207 57 213
rect 63 207 69 213
rect 75 207 81 213
rect 87 207 93 213
rect 99 207 105 213
rect 111 207 117 213
rect 123 207 129 213
rect 135 207 141 213
rect 147 207 153 213
rect 159 207 165 213
rect 171 207 177 213
rect 183 207 189 213
rect 195 207 201 213
rect 207 207 213 213
rect 219 207 225 213
rect 231 207 237 213
rect 243 207 249 213
rect 255 207 261 213
rect 267 207 273 213
rect 279 207 285 213
rect 291 207 297 213
rect 303 207 309 213
rect 315 207 321 213
rect 327 207 333 213
rect 339 207 345 213
rect 351 207 357 213
rect 363 207 369 213
rect 375 207 381 213
rect 387 207 393 213
rect 399 207 405 213
rect 411 207 417 213
rect 423 207 429 213
rect 435 207 441 213
rect 447 207 453 213
rect 459 207 465 213
rect 471 207 477 213
rect 483 207 489 213
rect 495 207 501 213
rect 507 207 513 213
rect 519 207 525 213
rect 531 207 537 213
rect 543 207 549 213
rect 555 207 561 213
rect 567 207 573 213
rect 579 207 585 213
rect 591 207 597 213
rect 603 207 609 213
rect 615 207 621 213
rect 627 207 633 213
rect 639 207 645 213
rect 651 207 657 213
rect 663 207 669 213
rect 675 207 681 213
rect 687 207 693 213
rect 699 207 705 213
rect 711 207 717 213
rect 723 207 729 213
rect 735 207 741 213
rect 747 207 753 213
rect 759 207 765 213
rect 771 207 777 213
rect 783 207 789 213
rect 795 207 801 213
rect 807 207 813 213
rect 819 207 825 213
rect 831 207 837 213
rect 843 207 849 213
rect 855 207 861 213
rect 867 207 873 213
rect 879 207 885 213
rect 891 207 897 213
rect 903 207 909 213
rect 915 207 921 213
rect 927 207 933 213
rect 939 207 945 213
rect 951 207 957 213
rect 963 207 969 213
rect 975 207 981 213
rect 987 207 993 213
rect 999 207 1005 213
rect 1011 207 1017 213
rect 1023 207 1029 213
rect 1035 207 1041 213
rect 1047 207 1053 213
rect 1059 207 1065 213
rect 1071 207 1077 213
rect 1083 207 1089 213
rect 1095 207 1101 213
rect 1107 207 1113 213
rect 1119 207 1125 213
rect 1131 207 1137 213
rect 1143 207 1149 213
rect 1155 207 1161 213
rect 1167 207 1173 213
rect 1179 207 1185 213
rect 1191 207 1197 213
rect 1203 207 1209 213
rect 1215 207 1221 213
rect 1227 207 1233 213
rect 1239 207 1245 213
rect 1251 207 1257 213
rect 1263 207 1269 213
rect 1275 207 1281 213
rect 1287 207 1293 213
rect 1299 207 1305 213
rect 1311 207 1317 213
rect 1323 207 1329 213
rect 1335 207 1341 213
rect 1347 207 1353 213
rect 1359 207 1365 213
rect 1371 207 1377 213
rect 1383 207 1389 213
rect 1395 207 1401 213
rect 1407 207 1413 213
rect 1419 207 1425 213
rect 1431 207 1437 213
rect 1443 207 1449 213
rect 1455 207 1461 213
rect 1467 207 1473 213
rect 1479 207 1485 213
rect 1491 207 1497 213
rect 1503 207 1509 213
rect 1515 207 1521 213
rect -45 87 -39 93
rect -33 87 -27 93
rect -21 87 -15 93
rect -9 87 -3 93
rect 3 87 9 93
rect 15 87 21 93
rect 27 87 33 93
rect 39 87 45 93
rect 51 87 57 93
rect 63 87 69 93
rect 75 87 81 93
rect 87 87 93 93
rect 99 87 105 93
rect 111 87 117 93
rect 123 87 129 93
rect 135 87 141 93
rect 147 87 153 93
rect 159 87 165 93
rect 171 87 177 93
rect 183 87 189 93
rect 195 87 201 93
rect 207 87 213 93
rect 219 87 225 93
rect 231 87 237 93
rect 243 87 249 93
rect 255 87 261 93
rect 267 87 273 93
rect 279 87 285 93
rect 291 87 297 93
rect 303 87 309 93
rect 315 87 321 93
rect 327 87 333 93
rect 339 87 345 93
rect 351 87 357 93
rect 363 87 369 93
rect 375 87 381 93
rect 387 87 393 93
rect 399 87 405 93
rect 411 87 417 93
rect 423 87 429 93
rect 435 87 441 93
rect 447 87 453 93
rect 459 87 465 93
rect 471 87 477 93
rect 483 87 489 93
rect 495 87 501 93
rect 507 87 513 93
rect 519 87 525 93
rect 531 87 537 93
rect 543 87 549 93
rect 555 87 561 93
rect 567 87 573 93
rect 579 87 585 93
rect 591 87 597 93
rect 603 87 609 93
rect 615 87 621 93
rect 627 87 633 93
rect 639 87 645 93
rect 651 87 657 93
rect 663 87 669 93
rect 675 87 681 93
rect 687 87 693 93
rect 699 87 705 93
rect 711 87 717 93
rect 723 87 729 93
rect 735 87 741 93
rect 747 87 753 93
rect 759 87 765 93
rect 771 87 777 93
rect 783 87 789 93
rect 795 87 801 93
rect 807 87 813 93
rect 819 87 825 93
rect 831 87 837 93
rect 843 87 849 93
rect 855 87 861 93
rect 867 87 873 93
rect 879 87 885 93
rect 891 87 897 93
rect 903 87 909 93
rect 915 87 921 93
rect 927 87 933 93
rect 939 87 945 93
rect 951 87 957 93
rect 963 87 969 93
rect 975 87 981 93
rect 987 87 993 93
rect 999 87 1005 93
rect 1011 87 1017 93
rect 1023 87 1029 93
rect 1035 87 1041 93
rect 1047 87 1053 93
rect 1059 87 1065 93
rect 1071 87 1077 93
rect 1083 87 1089 93
rect 1095 87 1101 93
rect 1107 87 1113 93
rect 1119 87 1125 93
rect 1131 87 1137 93
rect 1143 87 1149 93
rect 1155 87 1161 93
rect 1167 87 1173 93
rect 1179 87 1185 93
rect 1191 87 1197 93
rect 1203 87 1209 93
rect 1215 87 1221 93
rect 1227 87 1233 93
rect 1239 87 1245 93
rect 1251 87 1257 93
rect 1263 87 1269 93
rect 1275 87 1281 93
rect 1287 87 1293 93
rect 1299 87 1305 93
rect 1311 87 1317 93
rect 1323 87 1329 93
rect 1335 87 1341 93
rect 1347 87 1353 93
rect 1359 87 1365 93
rect 1371 87 1377 93
rect 1383 87 1389 93
rect 1395 87 1401 93
rect 1407 87 1413 93
rect 1419 87 1425 93
rect 1431 87 1437 93
rect 1443 87 1449 93
rect 1455 87 1461 93
rect 1467 87 1473 93
rect 1479 87 1485 93
rect 1491 87 1497 93
rect 1503 87 1509 93
rect 1515 87 1521 93
rect -45 -9 -39 -3
rect -33 -9 -27 -3
rect -21 -9 -15 -3
rect -9 -9 -3 -3
rect 3 -9 9 -3
rect 15 -9 21 -3
rect 27 -9 33 -3
rect 39 -9 45 -3
rect 51 -9 57 -3
rect 63 -9 69 -3
rect 75 -9 81 -3
rect 87 -9 93 -3
rect 99 -9 105 -3
rect 111 -9 117 -3
rect 123 -9 129 -3
rect 135 -9 141 -3
rect 147 -9 153 -3
rect 159 -9 165 -3
rect 171 -9 177 -3
rect 183 -9 189 -3
rect 195 -9 201 -3
rect 207 -9 213 -3
rect 219 -9 225 -3
rect 231 -9 237 -3
rect 243 -9 249 -3
rect 255 -9 261 -3
rect 267 -9 273 -3
rect 279 -9 285 -3
rect 291 -9 297 -3
rect 303 -9 309 -3
rect 315 -9 321 -3
rect 327 -9 333 -3
rect 339 -9 345 -3
rect 351 -9 357 -3
rect 363 -9 369 -3
rect 375 -9 381 -3
rect 387 -9 393 -3
rect 399 -9 405 -3
rect 411 -9 417 -3
rect 423 -9 429 -3
rect 435 -9 441 -3
rect 447 -9 453 -3
rect 459 -9 465 -3
rect 471 -9 477 -3
rect 483 -9 489 -3
rect 495 -9 501 -3
rect 507 -9 513 -3
rect 519 -9 525 -3
rect 531 -9 537 -3
rect 543 -9 549 -3
rect 555 -9 561 -3
rect 567 -9 573 -3
rect 579 -9 585 -3
rect 591 -9 597 -3
rect 603 -9 609 -3
rect 615 -9 621 -3
rect 627 -9 633 -3
rect 639 -9 645 -3
rect 651 -9 657 -3
rect 663 -9 669 -3
rect 675 -9 681 -3
rect 687 -9 693 -3
rect 699 -9 705 -3
rect 711 -9 717 -3
rect 723 -9 729 -3
rect 735 -9 741 -3
rect 747 -9 753 -3
rect 759 -9 765 -3
rect 771 -9 777 -3
rect 783 -9 789 -3
rect 795 -9 801 -3
rect 807 -9 813 -3
rect 819 -9 825 -3
rect 831 -9 837 -3
rect 843 -9 849 -3
rect 855 -9 861 -3
rect 867 -9 873 -3
rect 879 -9 885 -3
rect 891 -9 897 -3
rect 903 -9 909 -3
rect 915 -9 921 -3
rect 927 -9 933 -3
rect 939 -9 945 -3
rect 951 -9 957 -3
rect 963 -9 969 -3
rect 975 -9 981 -3
rect 987 -9 993 -3
rect 999 -9 1005 -3
rect 1011 -9 1017 -3
rect 1023 -9 1029 -3
rect 1035 -9 1041 -3
rect 1047 -9 1053 -3
rect 1059 -9 1065 -3
rect 1071 -9 1077 -3
rect 1083 -9 1089 -3
rect 1095 -9 1101 -3
rect 1107 -9 1113 -3
rect 1119 -9 1125 -3
rect 1131 -9 1137 -3
rect 1143 -9 1149 -3
rect 1155 -9 1161 -3
rect 1167 -9 1173 -3
rect 1179 -9 1185 -3
rect 1191 -9 1197 -3
rect 1203 -9 1209 -3
rect 1215 -9 1221 -3
rect 1227 -9 1233 -3
rect 1239 -9 1245 -3
rect 1251 -9 1257 -3
rect 1263 -9 1269 -3
rect 1275 -9 1281 -3
rect 1287 -9 1293 -3
rect 1299 -9 1305 -3
rect 1311 -9 1317 -3
rect 1323 -9 1329 -3
rect 1335 -9 1341 -3
rect 1347 -9 1353 -3
rect 1359 -9 1365 -3
rect 1371 -9 1377 -3
rect 1383 -9 1389 -3
rect 1395 -9 1401 -3
rect 1407 -9 1413 -3
rect 1419 -9 1425 -3
rect 1431 -9 1437 -3
rect 1443 -9 1449 -3
rect 1455 -9 1461 -3
rect 1467 -9 1473 -3
rect 1479 -9 1485 -3
rect 1491 -9 1497 -3
rect 1503 -9 1509 -3
rect 1515 -9 1521 -3
<< mvpsubdiffcont >>
rect -57 615 -51 621
rect -45 615 -39 621
rect -33 615 -27 621
rect -21 615 -15 621
rect -9 615 -3 621
rect 3 615 9 621
rect 15 615 21 621
rect 27 615 33 621
rect 39 615 45 621
rect 51 615 57 621
rect 63 615 69 621
rect 75 615 81 621
rect 87 615 93 621
rect 99 615 105 621
rect 111 615 117 621
rect 123 615 129 621
rect 135 615 141 621
rect 147 615 153 621
rect 159 615 165 621
rect 171 615 177 621
rect 183 615 189 621
rect 195 615 201 621
rect 207 615 213 621
rect 219 615 225 621
rect 231 615 237 621
rect 243 615 249 621
rect 255 615 261 621
rect 267 615 273 621
rect 279 615 285 621
rect 291 615 297 621
rect 303 615 309 621
rect 315 615 321 621
rect 327 615 333 621
rect 339 615 345 621
rect 351 615 357 621
rect 363 615 369 621
rect 375 615 381 621
rect 387 615 393 621
rect 399 615 405 621
rect 411 615 417 621
rect 423 615 429 621
rect 435 615 441 621
rect 447 615 453 621
rect 459 615 465 621
rect 471 615 477 621
rect 483 615 489 621
rect 495 615 501 621
rect 507 615 513 621
rect 519 615 525 621
rect 531 615 537 621
rect 543 615 549 621
rect 555 615 561 621
rect 567 615 573 621
rect 579 615 585 621
rect 591 615 597 621
rect 603 615 609 621
rect 615 615 621 621
rect 627 615 633 621
rect 639 615 645 621
rect 651 615 657 621
rect 663 615 669 621
rect 675 615 681 621
rect 687 615 693 621
rect 699 615 705 621
rect 711 615 717 621
rect 723 615 729 621
rect 735 615 741 621
rect 747 615 753 621
rect 759 615 765 621
rect 771 615 777 621
rect 783 615 789 621
rect 795 615 801 621
rect 807 615 813 621
rect 819 615 825 621
rect 831 615 837 621
rect 843 615 849 621
rect 855 615 861 621
rect 867 615 873 621
rect 879 615 885 621
rect 891 615 897 621
rect 903 615 909 621
rect 915 615 921 621
rect 927 615 933 621
rect 939 615 945 621
rect 951 615 957 621
rect 963 615 969 621
rect 975 615 981 621
rect 987 615 993 621
rect 999 615 1005 621
rect 1011 615 1017 621
rect 1023 615 1029 621
rect 1035 615 1041 621
rect 1047 615 1053 621
rect 1059 615 1065 621
rect 1071 615 1077 621
rect 1083 615 1089 621
rect 1095 615 1101 621
rect 1107 615 1113 621
rect 1119 615 1125 621
rect 1131 615 1137 621
rect 1143 615 1149 621
rect 1155 615 1161 621
rect 1167 615 1173 621
rect 1179 615 1185 621
rect 1191 615 1197 621
rect 1203 615 1209 621
rect 1215 615 1221 621
rect 1227 615 1233 621
rect 1239 615 1245 621
rect 1251 615 1257 621
rect 1263 615 1269 621
rect 1275 615 1281 621
rect 1287 615 1293 621
rect 1299 615 1305 621
rect 1311 615 1317 621
rect 1323 615 1329 621
rect 1335 615 1341 621
rect 1347 615 1353 621
rect 1359 615 1365 621
rect 1371 615 1377 621
rect 1383 615 1389 621
rect 1395 615 1401 621
rect 1407 615 1413 621
rect 1419 615 1425 621
rect 1431 615 1437 621
rect 1443 615 1449 621
rect 1455 615 1461 621
rect 1467 615 1473 621
rect 1479 615 1485 621
rect 1491 615 1497 621
rect 1503 615 1509 621
rect 1515 615 1521 621
rect 1527 615 1533 621
rect -57 603 -51 609
rect 1527 603 1533 609
rect -57 591 -51 597
rect -57 579 -51 585
rect -57 567 -51 573
rect -57 555 -51 561
rect -57 543 -51 549
rect -57 531 -51 537
rect -57 519 -51 525
rect -57 507 -51 513
rect -57 495 -51 501
rect -57 483 -51 489
rect -57 471 -51 477
rect -57 459 -51 465
rect -57 447 -51 453
rect -57 435 -51 441
rect -57 423 -51 429
rect -57 411 -51 417
rect -57 399 -51 405
rect -57 387 -51 393
rect -57 375 -51 381
rect -57 363 -51 369
rect -57 351 -51 357
rect 1527 591 1533 597
rect 1527 579 1533 585
rect 1527 567 1533 573
rect 1527 555 1533 561
rect 1527 543 1533 549
rect 1527 531 1533 537
rect 1527 519 1533 525
rect 1527 507 1533 513
rect 1527 495 1533 501
rect 1527 483 1533 489
rect 1527 471 1533 477
rect 1527 459 1533 465
rect 1527 447 1533 453
rect 1527 435 1533 441
rect 1527 423 1533 429
rect 1527 411 1533 417
rect 1527 399 1533 405
rect 1527 387 1533 393
rect 1527 375 1533 381
rect 1527 363 1533 369
rect 1527 351 1533 357
rect -57 339 -51 345
rect 1527 339 1533 345
rect -57 327 -51 333
rect -45 327 -39 333
rect -33 327 -27 333
rect -21 327 -15 333
rect -9 327 -3 333
rect 3 327 9 333
rect 15 327 21 333
rect 27 327 33 333
rect 39 327 45 333
rect 51 327 57 333
rect 63 327 69 333
rect 75 327 81 333
rect 87 327 93 333
rect 99 327 105 333
rect 111 327 117 333
rect 123 327 129 333
rect 135 327 141 333
rect 147 327 153 333
rect 159 327 165 333
rect 171 327 177 333
rect 183 327 189 333
rect 195 327 201 333
rect 207 327 213 333
rect 219 327 225 333
rect 231 327 237 333
rect 243 327 249 333
rect 255 327 261 333
rect 267 327 273 333
rect 279 327 285 333
rect 291 327 297 333
rect 303 327 309 333
rect 315 327 321 333
rect 327 327 333 333
rect 339 327 345 333
rect 351 327 357 333
rect 363 327 369 333
rect 375 327 381 333
rect 387 327 393 333
rect 399 327 405 333
rect 411 327 417 333
rect 423 327 429 333
rect 435 327 441 333
rect 447 327 453 333
rect 459 327 465 333
rect 471 327 477 333
rect 483 327 489 333
rect 495 327 501 333
rect 507 327 513 333
rect 519 327 525 333
rect 531 327 537 333
rect 543 327 549 333
rect 555 327 561 333
rect 567 327 573 333
rect 579 327 585 333
rect 591 327 597 333
rect 603 327 609 333
rect 615 327 621 333
rect 627 327 633 333
rect 639 327 645 333
rect 651 327 657 333
rect 663 327 669 333
rect 675 327 681 333
rect 687 327 693 333
rect 699 327 705 333
rect 711 327 717 333
rect 723 327 729 333
rect 735 327 741 333
rect 747 327 753 333
rect 759 327 765 333
rect 771 327 777 333
rect 783 327 789 333
rect 795 327 801 333
rect 807 327 813 333
rect 819 327 825 333
rect 831 327 837 333
rect 843 327 849 333
rect 855 327 861 333
rect 867 327 873 333
rect 879 327 885 333
rect 891 327 897 333
rect 903 327 909 333
rect 915 327 921 333
rect 927 327 933 333
rect 939 327 945 333
rect 951 327 957 333
rect 963 327 969 333
rect 975 327 981 333
rect 987 327 993 333
rect 999 327 1005 333
rect 1011 327 1017 333
rect 1023 327 1029 333
rect 1035 327 1041 333
rect 1047 327 1053 333
rect 1059 327 1065 333
rect 1071 327 1077 333
rect 1083 327 1089 333
rect 1095 327 1101 333
rect 1107 327 1113 333
rect 1119 327 1125 333
rect 1131 327 1137 333
rect 1143 327 1149 333
rect 1155 327 1161 333
rect 1167 327 1173 333
rect 1179 327 1185 333
rect 1191 327 1197 333
rect 1203 327 1209 333
rect 1215 327 1221 333
rect 1227 327 1233 333
rect 1239 327 1245 333
rect 1251 327 1257 333
rect 1263 327 1269 333
rect 1275 327 1281 333
rect 1287 327 1293 333
rect 1299 327 1305 333
rect 1311 327 1317 333
rect 1323 327 1329 333
rect 1335 327 1341 333
rect 1347 327 1353 333
rect 1359 327 1365 333
rect 1371 327 1377 333
rect 1383 327 1389 333
rect 1395 327 1401 333
rect 1407 327 1413 333
rect 1419 327 1425 333
rect 1431 327 1437 333
rect 1443 327 1449 333
rect 1455 327 1461 333
rect 1467 327 1473 333
rect 1479 327 1485 333
rect 1491 327 1497 333
rect 1503 327 1509 333
rect 1515 327 1521 333
rect 1527 327 1533 333
rect -57 315 -51 321
rect 1527 315 1533 321
rect -57 303 -51 309
rect -57 291 -51 297
rect 1527 303 1533 309
rect 1527 291 1533 297
rect -57 279 -51 285
rect -57 267 -51 273
rect -57 255 -51 261
rect 1527 279 1533 285
rect 1527 267 1533 273
rect 1527 255 1533 261
rect -57 243 -51 249
rect -57 231 -51 237
rect -57 219 -51 225
rect 1527 243 1533 249
rect 1527 231 1533 237
rect 1527 219 1533 225
rect -57 207 -51 213
rect 1527 207 1533 213
rect -57 195 -51 201
rect -57 183 -51 189
rect -57 171 -51 177
rect -57 159 -51 165
rect -57 147 -51 153
rect -57 135 -51 141
rect -57 123 -51 129
rect -57 111 -51 117
rect -57 99 -51 105
rect 1527 195 1533 201
rect 1527 183 1533 189
rect 1527 171 1533 177
rect 1527 159 1533 165
rect 1527 147 1533 153
rect 1527 135 1533 141
rect 1527 123 1533 129
rect 1527 111 1533 117
rect 1527 99 1533 105
rect -57 87 -51 93
rect 1527 87 1533 93
rect -57 75 -51 81
rect 1527 75 1533 81
rect -57 63 -51 69
rect -57 51 -51 57
rect 1527 63 1533 69
rect 1527 51 1533 57
rect -57 39 -51 45
rect -57 27 -51 33
rect -57 15 -51 21
rect 1527 39 1533 45
rect 1527 27 1533 33
rect 1527 15 1533 21
rect -57 3 -51 9
rect 1527 3 1533 9
rect -57 -9 -51 -3
rect 1527 -9 1533 -3
<< mvnsubdiffcont >>
rect -33 591 -27 597
rect -21 591 -15 597
rect -9 591 -3 597
rect 3 591 9 597
rect 15 591 21 597
rect 27 591 33 597
rect 39 591 45 597
rect 51 591 57 597
rect 63 591 69 597
rect 75 591 81 597
rect 87 591 93 597
rect 99 591 105 597
rect 111 591 117 597
rect 123 591 129 597
rect 135 591 141 597
rect 147 591 153 597
rect 159 591 165 597
rect 171 591 177 597
rect 183 591 189 597
rect 195 591 201 597
rect 207 591 213 597
rect 219 591 225 597
rect 231 591 237 597
rect 243 591 249 597
rect 255 591 261 597
rect 267 591 273 597
rect 279 591 285 597
rect 291 591 297 597
rect 303 591 309 597
rect 315 591 321 597
rect 327 591 333 597
rect 339 591 345 597
rect 351 591 357 597
rect 363 591 369 597
rect 375 591 381 597
rect 387 591 393 597
rect 399 591 405 597
rect 411 591 417 597
rect 423 591 429 597
rect 435 591 441 597
rect 447 591 453 597
rect 459 591 465 597
rect 471 591 477 597
rect 483 591 489 597
rect 495 591 501 597
rect 507 591 513 597
rect 519 591 525 597
rect 531 591 537 597
rect 543 591 549 597
rect 555 591 561 597
rect 567 591 573 597
rect 579 591 585 597
rect 591 591 597 597
rect 603 591 609 597
rect 615 591 621 597
rect 627 591 633 597
rect 639 591 645 597
rect 651 591 657 597
rect 663 591 669 597
rect 675 591 681 597
rect 687 591 693 597
rect 699 591 705 597
rect 711 591 717 597
rect 723 591 729 597
rect 735 591 741 597
rect 747 591 753 597
rect 759 591 765 597
rect 771 591 777 597
rect 783 591 789 597
rect 795 591 801 597
rect 807 591 813 597
rect 819 591 825 597
rect 831 591 837 597
rect 843 591 849 597
rect 855 591 861 597
rect 867 591 873 597
rect 879 591 885 597
rect 891 591 897 597
rect 903 591 909 597
rect 915 591 921 597
rect 927 591 933 597
rect 939 591 945 597
rect 951 591 957 597
rect 963 591 969 597
rect 975 591 981 597
rect 987 591 993 597
rect 999 591 1005 597
rect 1011 591 1017 597
rect 1023 591 1029 597
rect 1035 591 1041 597
rect 1047 591 1053 597
rect 1059 591 1065 597
rect 1071 591 1077 597
rect 1083 591 1089 597
rect 1095 591 1101 597
rect 1107 591 1113 597
rect 1119 591 1125 597
rect 1131 591 1137 597
rect 1143 591 1149 597
rect 1155 591 1161 597
rect 1167 591 1173 597
rect 1179 591 1185 597
rect 1191 591 1197 597
rect 1203 591 1209 597
rect 1215 591 1221 597
rect 1227 591 1233 597
rect 1239 591 1245 597
rect 1251 591 1257 597
rect 1263 591 1269 597
rect 1275 591 1281 597
rect 1287 591 1293 597
rect 1299 591 1305 597
rect 1311 591 1317 597
rect 1323 591 1329 597
rect 1335 591 1341 597
rect 1347 591 1353 597
rect 1359 591 1365 597
rect 1371 591 1377 597
rect 1383 591 1389 597
rect 1395 591 1401 597
rect 1407 591 1413 597
rect 1419 591 1425 597
rect 1431 591 1437 597
rect 1443 591 1449 597
rect 1455 591 1461 597
rect 1467 591 1473 597
rect 1479 591 1485 597
rect 1491 591 1497 597
rect 1503 591 1509 597
rect -33 579 -27 585
rect 1503 579 1509 585
rect -33 567 -27 573
rect -33 555 -27 561
rect -33 543 -27 549
rect 1503 567 1509 573
rect 1503 555 1509 561
rect 1503 543 1509 549
rect -33 531 -27 537
rect -33 519 -27 525
rect 1503 531 1509 537
rect 1503 519 1509 525
rect -33 507 -27 513
rect 1503 507 1509 513
rect -33 495 -27 501
rect -21 495 -15 501
rect -9 495 -3 501
rect 3 495 9 501
rect 15 495 21 501
rect 27 495 33 501
rect 39 495 45 501
rect 51 495 57 501
rect 63 495 69 501
rect 75 495 81 501
rect 87 495 93 501
rect 99 495 105 501
rect 111 495 117 501
rect 123 495 129 501
rect 135 495 141 501
rect 147 495 153 501
rect 159 495 165 501
rect 171 495 177 501
rect 183 495 189 501
rect 195 495 201 501
rect 207 495 213 501
rect 219 495 225 501
rect 231 495 237 501
rect 243 495 249 501
rect 255 495 261 501
rect 267 495 273 501
rect 279 495 285 501
rect 291 495 297 501
rect 303 495 309 501
rect 315 495 321 501
rect 327 495 333 501
rect 339 495 345 501
rect 351 495 357 501
rect 363 495 369 501
rect 375 495 381 501
rect 387 495 393 501
rect 399 495 405 501
rect 411 495 417 501
rect 423 495 429 501
rect 435 495 441 501
rect 447 495 453 501
rect 459 495 465 501
rect 471 495 477 501
rect 483 495 489 501
rect 495 495 501 501
rect 507 495 513 501
rect 519 495 525 501
rect 531 495 537 501
rect 543 495 549 501
rect 555 495 561 501
rect 567 495 573 501
rect 579 495 585 501
rect 591 495 597 501
rect 603 495 609 501
rect 615 495 621 501
rect 627 495 633 501
rect 639 495 645 501
rect 651 495 657 501
rect 663 495 669 501
rect 675 495 681 501
rect 687 495 693 501
rect 699 495 705 501
rect 711 495 717 501
rect 723 495 729 501
rect 735 495 741 501
rect 747 495 753 501
rect 759 495 765 501
rect 771 495 777 501
rect 783 495 789 501
rect 795 495 801 501
rect 807 495 813 501
rect 819 495 825 501
rect 831 495 837 501
rect 843 495 849 501
rect 855 495 861 501
rect 867 495 873 501
rect 879 495 885 501
rect 891 495 897 501
rect 903 495 909 501
rect 915 495 921 501
rect 927 495 933 501
rect 939 495 945 501
rect 951 495 957 501
rect 963 495 969 501
rect 975 495 981 501
rect 987 495 993 501
rect 999 495 1005 501
rect 1011 495 1017 501
rect 1023 495 1029 501
rect 1035 495 1041 501
rect 1047 495 1053 501
rect 1059 495 1065 501
rect 1071 495 1077 501
rect 1083 495 1089 501
rect 1095 495 1101 501
rect 1107 495 1113 501
rect 1119 495 1125 501
rect 1131 495 1137 501
rect 1143 495 1149 501
rect 1155 495 1161 501
rect 1167 495 1173 501
rect 1179 495 1185 501
rect 1191 495 1197 501
rect 1203 495 1209 501
rect 1215 495 1221 501
rect 1227 495 1233 501
rect 1239 495 1245 501
rect 1251 495 1257 501
rect 1263 495 1269 501
rect 1275 495 1281 501
rect 1287 495 1293 501
rect 1299 495 1305 501
rect 1311 495 1317 501
rect 1323 495 1329 501
rect 1335 495 1341 501
rect 1347 495 1353 501
rect 1359 495 1365 501
rect 1371 495 1377 501
rect 1383 495 1389 501
rect 1395 495 1401 501
rect 1407 495 1413 501
rect 1419 495 1425 501
rect 1431 495 1437 501
rect 1443 495 1449 501
rect 1455 495 1461 501
rect 1467 495 1473 501
rect 1479 495 1485 501
rect 1491 495 1497 501
rect 1503 495 1509 501
rect -33 483 -27 489
rect 1503 483 1509 489
rect -33 471 -27 477
rect -33 459 -27 465
rect -33 447 -27 453
rect 1503 471 1509 477
rect 1503 459 1509 465
rect 1503 447 1509 453
rect -33 435 -27 441
rect -33 423 -27 429
rect 1503 435 1509 441
rect 1503 423 1509 429
rect -33 411 -27 417
rect 1503 411 1509 417
rect -33 399 -27 405
rect -21 399 -15 405
rect -9 399 -3 405
rect 3 399 9 405
rect 15 399 21 405
rect 27 399 33 405
rect 39 399 45 405
rect 51 399 57 405
rect 63 399 69 405
rect 75 399 81 405
rect 87 399 93 405
rect 99 399 105 405
rect 111 399 117 405
rect 123 399 129 405
rect 135 399 141 405
rect 147 399 153 405
rect 159 399 165 405
rect 171 399 177 405
rect 183 399 189 405
rect 195 399 201 405
rect 207 399 213 405
rect 219 399 225 405
rect 231 399 237 405
rect 243 399 249 405
rect 255 399 261 405
rect 267 399 273 405
rect 279 399 285 405
rect 291 399 297 405
rect 303 399 309 405
rect 315 399 321 405
rect 327 399 333 405
rect 339 399 345 405
rect 351 399 357 405
rect 363 399 369 405
rect 375 399 381 405
rect 387 399 393 405
rect 399 399 405 405
rect 411 399 417 405
rect 423 399 429 405
rect 435 399 441 405
rect 447 399 453 405
rect 459 399 465 405
rect 471 399 477 405
rect 483 399 489 405
rect 495 399 501 405
rect 507 399 513 405
rect 519 399 525 405
rect 531 399 537 405
rect 543 399 549 405
rect 555 399 561 405
rect 567 399 573 405
rect 579 399 585 405
rect 591 399 597 405
rect 603 399 609 405
rect 615 399 621 405
rect 627 399 633 405
rect 639 399 645 405
rect 651 399 657 405
rect 663 399 669 405
rect 675 399 681 405
rect 687 399 693 405
rect 699 399 705 405
rect 711 399 717 405
rect 723 399 729 405
rect 735 399 741 405
rect 747 399 753 405
rect 759 399 765 405
rect 771 399 777 405
rect 783 399 789 405
rect 795 399 801 405
rect 807 399 813 405
rect 819 399 825 405
rect 831 399 837 405
rect 843 399 849 405
rect 855 399 861 405
rect 867 399 873 405
rect 879 399 885 405
rect 891 399 897 405
rect 903 399 909 405
rect 915 399 921 405
rect 927 399 933 405
rect 939 399 945 405
rect 951 399 957 405
rect 963 399 969 405
rect 975 399 981 405
rect 987 399 993 405
rect 999 399 1005 405
rect 1011 399 1017 405
rect 1023 399 1029 405
rect 1035 399 1041 405
rect 1047 399 1053 405
rect 1059 399 1065 405
rect 1071 399 1077 405
rect 1083 399 1089 405
rect 1095 399 1101 405
rect 1107 399 1113 405
rect 1119 399 1125 405
rect 1131 399 1137 405
rect 1143 399 1149 405
rect 1155 399 1161 405
rect 1167 399 1173 405
rect 1179 399 1185 405
rect 1191 399 1197 405
rect 1203 399 1209 405
rect 1215 399 1221 405
rect 1227 399 1233 405
rect 1239 399 1245 405
rect 1251 399 1257 405
rect 1263 399 1269 405
rect 1275 399 1281 405
rect 1287 399 1293 405
rect 1299 399 1305 405
rect 1311 399 1317 405
rect 1323 399 1329 405
rect 1335 399 1341 405
rect 1347 399 1353 405
rect 1359 399 1365 405
rect 1371 399 1377 405
rect 1383 399 1389 405
rect 1395 399 1401 405
rect 1407 399 1413 405
rect 1419 399 1425 405
rect 1431 399 1437 405
rect 1443 399 1449 405
rect 1455 399 1461 405
rect 1467 399 1473 405
rect 1479 399 1485 405
rect 1491 399 1497 405
rect 1503 399 1509 405
rect -33 387 -27 393
rect -33 375 -27 381
rect -33 363 -27 369
rect 1503 387 1509 393
rect 1503 375 1509 381
rect 1503 363 1509 369
rect -33 351 -27 357
rect -21 351 -15 357
rect -9 351 -3 357
rect 3 351 9 357
rect 15 351 21 357
rect 27 351 33 357
rect 39 351 45 357
rect 51 351 57 357
rect 63 351 69 357
rect 75 351 81 357
rect 87 351 93 357
rect 99 351 105 357
rect 111 351 117 357
rect 123 351 129 357
rect 135 351 141 357
rect 147 351 153 357
rect 159 351 165 357
rect 171 351 177 357
rect 183 351 189 357
rect 195 351 201 357
rect 207 351 213 357
rect 219 351 225 357
rect 231 351 237 357
rect 243 351 249 357
rect 255 351 261 357
rect 267 351 273 357
rect 279 351 285 357
rect 291 351 297 357
rect 303 351 309 357
rect 315 351 321 357
rect 327 351 333 357
rect 339 351 345 357
rect 351 351 357 357
rect 363 351 369 357
rect 375 351 381 357
rect 387 351 393 357
rect 399 351 405 357
rect 411 351 417 357
rect 423 351 429 357
rect 435 351 441 357
rect 447 351 453 357
rect 459 351 465 357
rect 471 351 477 357
rect 483 351 489 357
rect 495 351 501 357
rect 507 351 513 357
rect 519 351 525 357
rect 531 351 537 357
rect 543 351 549 357
rect 555 351 561 357
rect 567 351 573 357
rect 579 351 585 357
rect 591 351 597 357
rect 603 351 609 357
rect 615 351 621 357
rect 627 351 633 357
rect 639 351 645 357
rect 651 351 657 357
rect 663 351 669 357
rect 675 351 681 357
rect 687 351 693 357
rect 699 351 705 357
rect 711 351 717 357
rect 723 351 729 357
rect 735 351 741 357
rect 747 351 753 357
rect 759 351 765 357
rect 771 351 777 357
rect 783 351 789 357
rect 795 351 801 357
rect 807 351 813 357
rect 819 351 825 357
rect 831 351 837 357
rect 843 351 849 357
rect 855 351 861 357
rect 867 351 873 357
rect 879 351 885 357
rect 891 351 897 357
rect 903 351 909 357
rect 915 351 921 357
rect 927 351 933 357
rect 939 351 945 357
rect 951 351 957 357
rect 963 351 969 357
rect 975 351 981 357
rect 987 351 993 357
rect 999 351 1005 357
rect 1011 351 1017 357
rect 1023 351 1029 357
rect 1035 351 1041 357
rect 1047 351 1053 357
rect 1059 351 1065 357
rect 1071 351 1077 357
rect 1083 351 1089 357
rect 1095 351 1101 357
rect 1107 351 1113 357
rect 1119 351 1125 357
rect 1131 351 1137 357
rect 1143 351 1149 357
rect 1155 351 1161 357
rect 1167 351 1173 357
rect 1179 351 1185 357
rect 1191 351 1197 357
rect 1203 351 1209 357
rect 1215 351 1221 357
rect 1227 351 1233 357
rect 1239 351 1245 357
rect 1251 351 1257 357
rect 1263 351 1269 357
rect 1275 351 1281 357
rect 1287 351 1293 357
rect 1299 351 1305 357
rect 1311 351 1317 357
rect 1323 351 1329 357
rect 1335 351 1341 357
rect 1347 351 1353 357
rect 1359 351 1365 357
rect 1371 351 1377 357
rect 1383 351 1389 357
rect 1395 351 1401 357
rect 1407 351 1413 357
rect 1419 351 1425 357
rect 1431 351 1437 357
rect 1443 351 1449 357
rect 1455 351 1461 357
rect 1467 351 1473 357
rect 1479 351 1485 357
rect 1491 351 1497 357
rect 1503 351 1509 357
<< polysilicon >>
rect 0 576 12 582
rect 24 576 36 582
rect 48 576 60 582
rect 72 576 84 582
rect 96 576 108 582
rect 120 576 132 582
rect 144 576 156 582
rect 168 576 180 582
rect 216 576 228 582
rect 240 576 252 582
rect 264 576 276 582
rect 288 576 300 582
rect 312 576 324 582
rect 336 576 348 582
rect 360 576 372 582
rect 384 576 396 582
rect 432 576 444 582
rect 456 576 468 582
rect 480 576 492 582
rect 504 576 516 582
rect 528 576 540 582
rect 552 576 564 582
rect 576 576 588 582
rect 600 576 612 582
rect 648 576 660 582
rect 672 576 684 582
rect 696 576 708 582
rect 720 576 732 582
rect 744 576 756 582
rect 768 576 780 582
rect 792 576 804 582
rect 816 576 828 582
rect 864 576 876 582
rect 888 576 900 582
rect 912 576 924 582
rect 936 576 948 582
rect 960 576 972 582
rect 984 576 996 582
rect 1008 576 1020 582
rect 1032 576 1044 582
rect 1080 576 1092 582
rect 1104 576 1116 582
rect 1128 576 1140 582
rect 1152 576 1164 582
rect 1176 576 1188 582
rect 1200 576 1212 582
rect 1224 576 1236 582
rect 1248 576 1260 582
rect 1296 576 1308 582
rect 1320 576 1332 582
rect 1344 576 1356 582
rect 1368 576 1380 582
rect 1392 576 1404 582
rect 1416 576 1428 582
rect 1440 576 1452 582
rect 1464 576 1476 582
rect 0 528 12 540
rect 24 528 36 540
rect 0 525 36 528
rect 0 519 3 525
rect 9 519 15 525
rect 21 519 27 525
rect 33 519 36 525
rect 0 516 36 519
rect 48 528 60 540
rect 72 528 84 540
rect 48 525 84 528
rect 48 519 51 525
rect 57 519 63 525
rect 69 519 75 525
rect 81 519 84 525
rect 48 516 84 519
rect 96 528 108 540
rect 120 528 132 540
rect 96 525 132 528
rect 96 519 99 525
rect 105 519 111 525
rect 117 519 123 525
rect 129 519 132 525
rect 96 516 132 519
rect 144 528 156 540
rect 168 528 180 540
rect 144 525 180 528
rect 144 519 147 525
rect 153 519 159 525
rect 165 519 171 525
rect 177 519 180 525
rect 144 516 180 519
rect 216 528 228 540
rect 240 528 252 540
rect 216 525 252 528
rect 216 519 219 525
rect 225 519 231 525
rect 237 519 243 525
rect 249 519 252 525
rect 216 516 252 519
rect 264 528 276 540
rect 288 528 300 540
rect 264 525 300 528
rect 264 519 267 525
rect 273 519 279 525
rect 285 519 291 525
rect 297 519 300 525
rect 264 516 300 519
rect 312 528 324 540
rect 336 528 348 540
rect 312 525 348 528
rect 312 519 315 525
rect 321 519 327 525
rect 333 519 339 525
rect 345 519 348 525
rect 312 516 348 519
rect 360 528 372 540
rect 384 528 396 540
rect 360 525 396 528
rect 360 519 363 525
rect 369 519 375 525
rect 381 519 387 525
rect 393 519 396 525
rect 360 516 396 519
rect 432 528 444 540
rect 456 528 468 540
rect 432 525 468 528
rect 432 519 435 525
rect 441 519 447 525
rect 453 519 459 525
rect 465 519 468 525
rect 432 516 468 519
rect 480 528 492 540
rect 504 528 516 540
rect 480 525 516 528
rect 480 519 483 525
rect 489 519 495 525
rect 501 519 507 525
rect 513 519 516 525
rect 480 516 516 519
rect 528 528 540 540
rect 552 528 564 540
rect 528 525 564 528
rect 528 519 531 525
rect 537 519 543 525
rect 549 519 555 525
rect 561 519 564 525
rect 528 516 564 519
rect 576 528 588 540
rect 600 528 612 540
rect 576 525 612 528
rect 576 519 579 525
rect 585 519 591 525
rect 597 519 603 525
rect 609 519 612 525
rect 576 516 612 519
rect 648 528 660 540
rect 672 528 684 540
rect 648 525 684 528
rect 648 519 651 525
rect 657 519 663 525
rect 669 519 675 525
rect 681 519 684 525
rect 648 516 684 519
rect 696 528 708 540
rect 720 528 732 540
rect 696 525 732 528
rect 696 519 699 525
rect 705 519 711 525
rect 717 519 723 525
rect 729 519 732 525
rect 696 516 732 519
rect 744 528 756 540
rect 768 528 780 540
rect 744 525 780 528
rect 744 519 747 525
rect 753 519 759 525
rect 765 519 771 525
rect 777 519 780 525
rect 744 516 780 519
rect 792 528 804 540
rect 816 528 828 540
rect 792 525 828 528
rect 792 519 795 525
rect 801 519 807 525
rect 813 519 819 525
rect 825 519 828 525
rect 792 516 828 519
rect 864 528 876 540
rect 888 528 900 540
rect 912 528 924 540
rect 936 528 948 540
rect 864 525 948 528
rect 864 519 867 525
rect 873 519 879 525
rect 885 519 891 525
rect 897 519 903 525
rect 909 519 915 525
rect 921 519 927 525
rect 933 519 939 525
rect 945 519 948 525
rect 864 516 948 519
rect 960 528 972 540
rect 984 528 996 540
rect 960 525 996 528
rect 960 519 963 525
rect 969 519 975 525
rect 981 519 987 525
rect 993 519 996 525
rect 960 516 996 519
rect 1008 528 1020 540
rect 1032 528 1044 540
rect 1008 525 1044 528
rect 1008 519 1011 525
rect 1017 519 1023 525
rect 1029 519 1035 525
rect 1041 519 1044 525
rect 1008 516 1044 519
rect 1080 528 1092 540
rect 1104 528 1116 540
rect 1080 525 1116 528
rect 1080 519 1083 525
rect 1089 519 1095 525
rect 1101 519 1107 525
rect 1113 519 1116 525
rect 1080 516 1116 519
rect 1128 528 1140 540
rect 1152 528 1164 540
rect 1128 525 1164 528
rect 1128 519 1131 525
rect 1137 519 1143 525
rect 1149 519 1155 525
rect 1161 519 1164 525
rect 1128 516 1164 519
rect 1176 528 1188 540
rect 1200 528 1212 540
rect 1176 525 1212 528
rect 1176 519 1179 525
rect 1185 519 1191 525
rect 1197 519 1203 525
rect 1209 519 1212 525
rect 1176 516 1212 519
rect 1224 528 1236 540
rect 1248 528 1260 540
rect 1224 525 1260 528
rect 1224 519 1227 525
rect 1233 519 1239 525
rect 1245 519 1251 525
rect 1257 519 1260 525
rect 1224 516 1260 519
rect 1296 528 1308 540
rect 1320 528 1332 540
rect 1296 525 1332 528
rect 1296 519 1299 525
rect 1305 519 1311 525
rect 1317 519 1323 525
rect 1329 519 1332 525
rect 1296 516 1332 519
rect 1344 528 1356 540
rect 1368 528 1380 540
rect 1344 525 1380 528
rect 1344 519 1347 525
rect 1353 519 1359 525
rect 1365 519 1371 525
rect 1377 519 1380 525
rect 1344 516 1380 519
rect 1392 528 1404 540
rect 1416 528 1428 540
rect 1392 525 1428 528
rect 1392 519 1395 525
rect 1401 519 1407 525
rect 1413 519 1419 525
rect 1425 519 1428 525
rect 1392 516 1428 519
rect 1440 528 1452 540
rect 1464 528 1476 540
rect 1440 525 1476 528
rect 1440 519 1443 525
rect 1449 519 1455 525
rect 1461 519 1467 525
rect 1473 519 1476 525
rect 1440 516 1476 519
rect 0 480 12 486
rect 24 480 36 486
rect 48 480 60 486
rect 72 480 84 486
rect 96 480 108 486
rect 120 480 132 486
rect 144 480 156 486
rect 168 480 180 486
rect 216 480 228 486
rect 240 480 252 486
rect 264 480 276 486
rect 288 480 300 486
rect 312 480 324 486
rect 336 480 348 486
rect 360 480 372 486
rect 384 480 396 486
rect 432 480 444 486
rect 456 480 468 486
rect 480 480 492 486
rect 504 480 516 486
rect 528 480 540 486
rect 552 480 564 486
rect 576 480 588 486
rect 600 480 612 486
rect 648 480 660 486
rect 672 480 684 486
rect 696 480 708 486
rect 720 480 732 486
rect 744 480 756 486
rect 768 480 780 486
rect 792 480 804 486
rect 816 480 828 486
rect 864 480 876 486
rect 888 480 900 486
rect 912 480 924 486
rect 936 480 948 486
rect 960 480 972 486
rect 984 480 996 486
rect 1008 480 1020 486
rect 1032 480 1044 486
rect 1080 480 1092 486
rect 1104 480 1116 486
rect 1128 480 1140 486
rect 1152 480 1164 486
rect 1176 480 1188 486
rect 1200 480 1212 486
rect 1224 480 1236 486
rect 1248 480 1260 486
rect 1296 480 1308 486
rect 1320 480 1332 486
rect 1344 480 1356 486
rect 1368 480 1380 486
rect 1392 480 1404 486
rect 1416 480 1428 486
rect 1440 480 1452 486
rect 1464 480 1476 486
rect 0 432 12 444
rect 24 432 36 444
rect 0 429 36 432
rect 0 423 3 429
rect 9 423 15 429
rect 21 423 27 429
rect 33 423 36 429
rect 0 420 36 423
rect 48 432 60 444
rect 72 432 84 444
rect 48 429 84 432
rect 48 423 51 429
rect 57 423 63 429
rect 69 423 75 429
rect 81 423 84 429
rect 48 420 84 423
rect 96 432 108 444
rect 120 432 132 444
rect 96 429 132 432
rect 96 423 99 429
rect 105 423 111 429
rect 117 423 123 429
rect 129 423 132 429
rect 96 420 132 423
rect 144 432 156 444
rect 168 432 180 444
rect 144 429 180 432
rect 144 423 147 429
rect 153 423 159 429
rect 165 423 171 429
rect 177 423 180 429
rect 144 420 180 423
rect 216 432 228 444
rect 240 432 252 444
rect 216 429 252 432
rect 216 423 219 429
rect 225 423 231 429
rect 237 423 243 429
rect 249 423 252 429
rect 216 420 252 423
rect 264 432 276 444
rect 288 432 300 444
rect 264 429 300 432
rect 264 423 267 429
rect 273 423 279 429
rect 285 423 291 429
rect 297 423 300 429
rect 264 420 300 423
rect 312 432 324 444
rect 336 432 348 444
rect 312 429 348 432
rect 312 423 315 429
rect 321 423 327 429
rect 333 423 339 429
rect 345 423 348 429
rect 312 420 348 423
rect 360 432 372 444
rect 384 432 396 444
rect 360 429 396 432
rect 360 423 363 429
rect 369 423 375 429
rect 381 423 387 429
rect 393 423 396 429
rect 360 420 396 423
rect 432 432 444 444
rect 456 432 468 444
rect 432 429 468 432
rect 432 423 435 429
rect 441 423 447 429
rect 453 423 459 429
rect 465 423 468 429
rect 432 420 468 423
rect 480 432 492 444
rect 504 432 516 444
rect 480 429 516 432
rect 480 423 483 429
rect 489 423 495 429
rect 501 423 507 429
rect 513 423 516 429
rect 480 420 516 423
rect 528 432 540 444
rect 552 432 564 444
rect 528 429 564 432
rect 528 423 531 429
rect 537 423 543 429
rect 549 423 555 429
rect 561 423 564 429
rect 528 420 564 423
rect 576 432 588 444
rect 600 432 612 444
rect 576 429 612 432
rect 576 423 579 429
rect 585 423 591 429
rect 597 423 603 429
rect 609 423 612 429
rect 576 420 612 423
rect 648 432 660 444
rect 672 432 684 444
rect 648 429 684 432
rect 648 423 651 429
rect 657 423 663 429
rect 669 423 675 429
rect 681 423 684 429
rect 648 420 684 423
rect 696 432 708 444
rect 720 432 732 444
rect 696 429 732 432
rect 696 423 699 429
rect 705 423 711 429
rect 717 423 723 429
rect 729 423 732 429
rect 696 420 732 423
rect 744 432 756 444
rect 768 432 780 444
rect 744 429 780 432
rect 744 423 747 429
rect 753 423 759 429
rect 765 423 771 429
rect 777 423 780 429
rect 744 420 780 423
rect 792 432 804 444
rect 816 432 828 444
rect 792 429 828 432
rect 792 423 795 429
rect 801 423 807 429
rect 813 423 819 429
rect 825 423 828 429
rect 792 420 828 423
rect 864 432 876 444
rect 888 432 900 444
rect 912 432 924 444
rect 936 432 948 444
rect 864 429 948 432
rect 864 423 867 429
rect 873 423 879 429
rect 885 423 891 429
rect 897 423 903 429
rect 909 423 915 429
rect 921 423 927 429
rect 933 423 939 429
rect 945 423 948 429
rect 864 420 948 423
rect 960 432 972 444
rect 984 432 996 444
rect 960 429 996 432
rect 960 423 963 429
rect 969 423 975 429
rect 981 423 987 429
rect 993 423 996 429
rect 960 420 996 423
rect 1008 432 1020 444
rect 1032 432 1044 444
rect 1008 429 1044 432
rect 1008 423 1011 429
rect 1017 423 1023 429
rect 1029 423 1035 429
rect 1041 423 1044 429
rect 1008 420 1044 423
rect 1080 432 1092 444
rect 1104 432 1116 444
rect 1080 429 1116 432
rect 1080 423 1083 429
rect 1089 423 1095 429
rect 1101 423 1107 429
rect 1113 423 1116 429
rect 1080 420 1116 423
rect 1128 432 1140 444
rect 1152 432 1164 444
rect 1128 429 1164 432
rect 1128 423 1131 429
rect 1137 423 1143 429
rect 1149 423 1155 429
rect 1161 423 1164 429
rect 1128 420 1164 423
rect 1176 432 1188 444
rect 1200 432 1212 444
rect 1176 429 1212 432
rect 1176 423 1179 429
rect 1185 423 1191 429
rect 1197 423 1203 429
rect 1209 423 1212 429
rect 1176 420 1212 423
rect 1224 432 1236 444
rect 1248 432 1260 444
rect 1224 429 1260 432
rect 1224 423 1227 429
rect 1233 423 1239 429
rect 1245 423 1251 429
rect 1257 423 1260 429
rect 1224 420 1260 423
rect 1296 432 1308 444
rect 1320 432 1332 444
rect 1296 429 1332 432
rect 1296 423 1299 429
rect 1305 423 1311 429
rect 1317 423 1323 429
rect 1329 423 1332 429
rect 1296 420 1332 423
rect 1344 432 1356 444
rect 1368 432 1380 444
rect 1344 429 1380 432
rect 1344 423 1347 429
rect 1353 423 1359 429
rect 1365 423 1371 429
rect 1377 423 1380 429
rect 1344 420 1380 423
rect 1392 432 1404 444
rect 1416 432 1428 444
rect 1392 429 1428 432
rect 1392 423 1395 429
rect 1401 423 1407 429
rect 1413 423 1419 429
rect 1425 423 1428 429
rect 1392 420 1428 423
rect 1440 432 1452 444
rect 1464 432 1476 444
rect 1440 429 1476 432
rect 1440 423 1443 429
rect 1449 423 1455 429
rect 1461 423 1467 429
rect 1473 423 1476 429
rect 1440 420 1476 423
rect 0 309 36 312
rect 0 303 3 309
rect 9 303 15 309
rect 21 303 27 309
rect 33 303 36 309
rect 0 300 36 303
rect 0 288 12 300
rect 24 288 36 300
rect 48 309 84 312
rect 48 303 51 309
rect 57 303 63 309
rect 69 303 75 309
rect 81 303 84 309
rect 48 300 84 303
rect 48 288 60 300
rect 72 288 84 300
rect 96 309 132 312
rect 96 303 99 309
rect 105 303 111 309
rect 117 303 123 309
rect 129 303 132 309
rect 96 300 132 303
rect 96 288 108 300
rect 120 288 132 300
rect 144 309 180 312
rect 144 303 147 309
rect 153 303 159 309
rect 165 303 171 309
rect 177 303 180 309
rect 144 300 180 303
rect 144 288 156 300
rect 168 288 180 300
rect 216 309 252 312
rect 216 303 219 309
rect 225 303 231 309
rect 237 303 243 309
rect 249 303 252 309
rect 216 300 252 303
rect 216 288 228 300
rect 240 288 252 300
rect 264 309 300 312
rect 264 303 267 309
rect 273 303 279 309
rect 285 303 291 309
rect 297 303 300 309
rect 264 300 300 303
rect 264 288 276 300
rect 288 288 300 300
rect 312 309 348 312
rect 312 303 315 309
rect 321 303 327 309
rect 333 303 339 309
rect 345 303 348 309
rect 312 300 348 303
rect 312 288 324 300
rect 336 288 348 300
rect 360 309 396 312
rect 360 303 363 309
rect 369 303 375 309
rect 381 303 387 309
rect 393 303 396 309
rect 360 300 396 303
rect 360 288 372 300
rect 384 288 396 300
rect 432 309 468 312
rect 432 303 435 309
rect 441 303 447 309
rect 453 303 459 309
rect 465 303 468 309
rect 432 300 468 303
rect 432 288 444 300
rect 456 288 468 300
rect 480 309 516 312
rect 480 303 483 309
rect 489 303 495 309
rect 501 303 507 309
rect 513 303 516 309
rect 480 300 516 303
rect 480 288 492 300
rect 504 288 516 300
rect 528 309 564 312
rect 528 303 531 309
rect 537 303 543 309
rect 549 303 555 309
rect 561 303 564 309
rect 528 300 564 303
rect 528 288 540 300
rect 552 288 564 300
rect 576 309 612 312
rect 576 303 579 309
rect 585 303 591 309
rect 597 303 603 309
rect 609 303 612 309
rect 576 300 612 303
rect 576 288 588 300
rect 600 288 612 300
rect 648 309 684 312
rect 648 303 651 309
rect 657 303 663 309
rect 669 303 675 309
rect 681 303 684 309
rect 648 300 684 303
rect 648 288 660 300
rect 672 288 684 300
rect 696 309 732 312
rect 696 303 699 309
rect 705 303 711 309
rect 717 303 723 309
rect 729 303 732 309
rect 696 300 732 303
rect 696 288 708 300
rect 720 288 732 300
rect 744 309 780 312
rect 744 303 747 309
rect 753 303 759 309
rect 765 303 771 309
rect 777 303 780 309
rect 744 300 780 303
rect 744 288 756 300
rect 768 288 780 300
rect 792 309 828 312
rect 792 303 795 309
rect 801 303 807 309
rect 813 303 819 309
rect 825 303 828 309
rect 792 300 828 303
rect 792 288 804 300
rect 816 288 828 300
rect 864 309 876 312
rect 864 303 867 309
rect 873 303 876 309
rect 864 288 876 303
rect 912 309 948 312
rect 912 303 915 309
rect 921 303 927 309
rect 933 303 939 309
rect 945 303 948 309
rect 912 300 948 303
rect 912 288 924 300
rect 936 288 948 300
rect 960 309 996 312
rect 960 303 963 309
rect 969 303 975 309
rect 981 303 987 309
rect 993 303 996 309
rect 960 300 996 303
rect 960 288 972 300
rect 984 288 996 300
rect 1008 309 1044 312
rect 1008 303 1011 309
rect 1017 303 1023 309
rect 1029 303 1035 309
rect 1041 303 1044 309
rect 1008 300 1044 303
rect 1008 288 1020 300
rect 1032 288 1044 300
rect 1080 309 1116 312
rect 1080 303 1083 309
rect 1089 303 1095 309
rect 1101 303 1107 309
rect 1113 303 1116 309
rect 1080 300 1116 303
rect 1080 288 1092 300
rect 1104 288 1116 300
rect 1128 309 1164 312
rect 1128 303 1131 309
rect 1137 303 1143 309
rect 1149 303 1155 309
rect 1161 303 1164 309
rect 1128 300 1164 303
rect 1128 288 1140 300
rect 1152 288 1164 300
rect 1176 309 1212 312
rect 1176 303 1179 309
rect 1185 303 1191 309
rect 1197 303 1203 309
rect 1209 303 1212 309
rect 1176 300 1212 303
rect 1176 288 1188 300
rect 1200 288 1212 300
rect 1224 309 1260 312
rect 1224 303 1227 309
rect 1233 303 1239 309
rect 1245 303 1251 309
rect 1257 303 1260 309
rect 1224 300 1260 303
rect 1224 288 1236 300
rect 1248 288 1260 300
rect 1296 309 1332 312
rect 1296 303 1299 309
rect 1305 303 1311 309
rect 1317 303 1323 309
rect 1329 303 1332 309
rect 1296 300 1332 303
rect 1296 288 1308 300
rect 1320 288 1332 300
rect 1344 309 1380 312
rect 1344 303 1347 309
rect 1353 303 1359 309
rect 1365 303 1371 309
rect 1377 303 1380 309
rect 1344 300 1380 303
rect 1344 288 1356 300
rect 1368 288 1380 300
rect 1392 309 1428 312
rect 1392 303 1395 309
rect 1401 303 1407 309
rect 1413 303 1419 309
rect 1425 303 1428 309
rect 1392 300 1428 303
rect 1392 288 1404 300
rect 1416 288 1428 300
rect 1440 309 1476 312
rect 1440 303 1443 309
rect 1449 303 1455 309
rect 1461 303 1467 309
rect 1473 303 1476 309
rect 1440 300 1476 303
rect 1440 288 1452 300
rect 1464 288 1476 300
rect 0 246 12 252
rect 24 246 36 252
rect 48 246 60 252
rect 72 246 84 252
rect 96 246 108 252
rect 120 246 132 252
rect 144 246 156 252
rect 168 246 180 252
rect 216 246 228 252
rect 240 246 252 252
rect 264 246 276 252
rect 288 246 300 252
rect 312 246 324 252
rect 336 246 348 252
rect 360 246 372 252
rect 384 246 396 252
rect 432 246 444 252
rect 456 246 468 252
rect 480 246 492 252
rect 504 246 516 252
rect 528 246 540 252
rect 552 246 564 252
rect 576 246 588 252
rect 600 246 612 252
rect 648 246 660 252
rect 672 246 684 252
rect 696 246 708 252
rect 720 246 732 252
rect 744 246 756 252
rect 768 246 780 252
rect 792 246 804 252
rect 816 246 828 252
rect 864 246 876 252
rect 912 246 924 252
rect 936 246 948 252
rect 960 246 972 252
rect 984 246 996 252
rect 1008 246 1020 252
rect 1032 246 1044 252
rect 1080 246 1092 252
rect 1104 246 1116 252
rect 1128 246 1140 252
rect 1152 246 1164 252
rect 1176 246 1188 252
rect 1200 246 1212 252
rect 1224 246 1236 252
rect 1248 246 1260 252
rect 1296 246 1308 252
rect 1320 246 1332 252
rect 1344 246 1356 252
rect 1368 246 1380 252
rect 1392 246 1404 252
rect 1416 246 1428 252
rect 1440 246 1452 252
rect 1464 246 1476 252
rect 0 69 36 72
rect 0 63 3 69
rect 9 63 15 69
rect 21 63 27 69
rect 33 63 36 69
rect 0 60 36 63
rect 0 48 12 60
rect 24 48 36 60
rect 48 69 84 72
rect 48 63 51 69
rect 57 63 63 69
rect 69 63 75 69
rect 81 63 84 69
rect 48 60 84 63
rect 48 48 60 60
rect 72 48 84 60
rect 96 69 132 72
rect 96 63 99 69
rect 105 63 111 69
rect 117 63 123 69
rect 129 63 132 69
rect 96 60 132 63
rect 96 48 108 60
rect 120 48 132 60
rect 144 69 180 72
rect 144 63 147 69
rect 153 63 159 69
rect 165 63 171 69
rect 177 63 180 69
rect 144 60 180 63
rect 144 48 156 60
rect 168 48 180 60
rect 216 69 252 72
rect 216 63 219 69
rect 225 63 231 69
rect 237 63 243 69
rect 249 63 252 69
rect 216 60 252 63
rect 216 48 228 60
rect 240 48 252 60
rect 264 69 300 72
rect 264 63 267 69
rect 273 63 279 69
rect 285 63 291 69
rect 297 63 300 69
rect 264 60 300 63
rect 264 48 276 60
rect 288 48 300 60
rect 312 69 348 72
rect 312 63 315 69
rect 321 63 327 69
rect 333 63 339 69
rect 345 63 348 69
rect 312 60 348 63
rect 312 48 324 60
rect 336 48 348 60
rect 360 69 396 72
rect 360 63 363 69
rect 369 63 375 69
rect 381 63 387 69
rect 393 63 396 69
rect 360 60 396 63
rect 360 48 372 60
rect 384 48 396 60
rect 432 69 468 72
rect 432 63 435 69
rect 441 63 447 69
rect 453 63 459 69
rect 465 63 468 69
rect 432 60 468 63
rect 432 48 444 60
rect 456 48 468 60
rect 480 69 516 72
rect 480 63 483 69
rect 489 63 495 69
rect 501 63 507 69
rect 513 63 516 69
rect 480 60 516 63
rect 480 48 492 60
rect 504 48 516 60
rect 528 69 564 72
rect 528 63 531 69
rect 537 63 543 69
rect 549 63 555 69
rect 561 63 564 69
rect 528 60 564 63
rect 528 48 540 60
rect 552 48 564 60
rect 576 69 612 72
rect 576 63 579 69
rect 585 63 591 69
rect 597 63 603 69
rect 609 63 612 69
rect 576 60 612 63
rect 576 48 588 60
rect 600 48 612 60
rect 648 69 684 72
rect 648 63 651 69
rect 657 63 663 69
rect 669 63 675 69
rect 681 63 684 69
rect 648 60 684 63
rect 648 48 660 60
rect 672 48 684 60
rect 696 69 732 72
rect 696 63 699 69
rect 705 63 711 69
rect 717 63 723 69
rect 729 63 732 69
rect 696 60 732 63
rect 696 48 708 60
rect 720 48 732 60
rect 744 69 780 72
rect 744 63 747 69
rect 753 63 759 69
rect 765 63 771 69
rect 777 63 780 69
rect 744 60 780 63
rect 744 48 756 60
rect 768 48 780 60
rect 792 69 828 72
rect 792 63 795 69
rect 801 63 807 69
rect 813 63 819 69
rect 825 63 828 69
rect 792 60 828 63
rect 792 48 804 60
rect 816 48 828 60
rect 864 69 900 72
rect 864 63 867 69
rect 873 63 879 69
rect 885 63 891 69
rect 897 63 900 69
rect 864 60 900 63
rect 864 48 876 60
rect 888 48 900 60
rect 912 69 948 72
rect 912 63 915 69
rect 921 63 927 69
rect 933 63 939 69
rect 945 63 948 69
rect 912 60 948 63
rect 912 48 924 60
rect 936 48 948 60
rect 960 69 996 72
rect 960 63 963 69
rect 969 63 975 69
rect 981 63 987 69
rect 993 63 996 69
rect 960 60 996 63
rect 960 48 972 60
rect 984 48 996 60
rect 1008 69 1044 72
rect 1008 63 1011 69
rect 1017 63 1023 69
rect 1029 63 1035 69
rect 1041 63 1044 69
rect 1008 60 1044 63
rect 1008 48 1020 60
rect 1032 48 1044 60
rect 1080 69 1116 72
rect 1080 63 1083 69
rect 1089 63 1095 69
rect 1101 63 1107 69
rect 1113 63 1116 69
rect 1080 60 1116 63
rect 1080 48 1092 60
rect 1104 48 1116 60
rect 1128 69 1164 72
rect 1128 63 1131 69
rect 1137 63 1143 69
rect 1149 63 1155 69
rect 1161 63 1164 69
rect 1128 60 1164 63
rect 1128 48 1140 60
rect 1152 48 1164 60
rect 1176 69 1212 72
rect 1176 63 1179 69
rect 1185 63 1191 69
rect 1197 63 1203 69
rect 1209 63 1212 69
rect 1176 60 1212 63
rect 1176 48 1188 60
rect 1200 48 1212 60
rect 1224 69 1260 72
rect 1224 63 1227 69
rect 1233 63 1239 69
rect 1245 63 1251 69
rect 1257 63 1260 69
rect 1224 60 1260 63
rect 1224 48 1236 60
rect 1248 48 1260 60
rect 1296 69 1332 72
rect 1296 63 1299 69
rect 1305 63 1311 69
rect 1317 63 1323 69
rect 1329 63 1332 69
rect 1296 60 1332 63
rect 1296 48 1308 60
rect 1320 48 1332 60
rect 1344 69 1380 72
rect 1344 63 1347 69
rect 1353 63 1359 69
rect 1365 63 1371 69
rect 1377 63 1380 69
rect 1344 60 1380 63
rect 1344 48 1356 60
rect 1368 48 1380 60
rect 1392 69 1428 72
rect 1392 63 1395 69
rect 1401 63 1407 69
rect 1413 63 1419 69
rect 1425 63 1428 69
rect 1392 60 1428 63
rect 1392 48 1404 60
rect 1416 48 1428 60
rect 1440 69 1476 72
rect 1440 63 1443 69
rect 1449 63 1455 69
rect 1461 63 1467 69
rect 1473 63 1476 69
rect 1440 60 1476 63
rect 1440 48 1452 60
rect 1464 48 1476 60
rect 0 6 12 12
rect 24 6 36 12
rect 48 6 60 12
rect 72 6 84 12
rect 96 6 108 12
rect 120 6 132 12
rect 144 6 156 12
rect 168 6 180 12
rect 216 6 228 12
rect 240 6 252 12
rect 264 6 276 12
rect 288 6 300 12
rect 312 6 324 12
rect 336 6 348 12
rect 360 6 372 12
rect 384 6 396 12
rect 432 6 444 12
rect 456 6 468 12
rect 480 6 492 12
rect 504 6 516 12
rect 528 6 540 12
rect 552 6 564 12
rect 576 6 588 12
rect 600 6 612 12
rect 648 6 660 12
rect 672 6 684 12
rect 696 6 708 12
rect 720 6 732 12
rect 744 6 756 12
rect 768 6 780 12
rect 792 6 804 12
rect 816 6 828 12
rect 864 6 876 12
rect 888 6 900 12
rect 912 6 924 12
rect 936 6 948 12
rect 960 6 972 12
rect 984 6 996 12
rect 1008 6 1020 12
rect 1032 6 1044 12
rect 1080 6 1092 12
rect 1104 6 1116 12
rect 1128 6 1140 12
rect 1152 6 1164 12
rect 1176 6 1188 12
rect 1200 6 1212 12
rect 1224 6 1236 12
rect 1248 6 1260 12
rect 1296 6 1308 12
rect 1320 6 1332 12
rect 1344 6 1356 12
rect 1368 6 1380 12
rect 1392 6 1404 12
rect 1416 6 1428 12
rect 1440 6 1452 12
rect 1464 6 1476 12
<< polycontact >>
rect 3 519 9 525
rect 15 519 21 525
rect 27 519 33 525
rect 51 519 57 525
rect 63 519 69 525
rect 75 519 81 525
rect 99 519 105 525
rect 111 519 117 525
rect 123 519 129 525
rect 147 519 153 525
rect 159 519 165 525
rect 171 519 177 525
rect 219 519 225 525
rect 231 519 237 525
rect 243 519 249 525
rect 267 519 273 525
rect 279 519 285 525
rect 291 519 297 525
rect 315 519 321 525
rect 327 519 333 525
rect 339 519 345 525
rect 363 519 369 525
rect 375 519 381 525
rect 387 519 393 525
rect 435 519 441 525
rect 447 519 453 525
rect 459 519 465 525
rect 483 519 489 525
rect 495 519 501 525
rect 507 519 513 525
rect 531 519 537 525
rect 543 519 549 525
rect 555 519 561 525
rect 579 519 585 525
rect 591 519 597 525
rect 603 519 609 525
rect 651 519 657 525
rect 663 519 669 525
rect 675 519 681 525
rect 699 519 705 525
rect 711 519 717 525
rect 723 519 729 525
rect 747 519 753 525
rect 759 519 765 525
rect 771 519 777 525
rect 795 519 801 525
rect 807 519 813 525
rect 819 519 825 525
rect 867 519 873 525
rect 879 519 885 525
rect 891 519 897 525
rect 903 519 909 525
rect 915 519 921 525
rect 927 519 933 525
rect 939 519 945 525
rect 963 519 969 525
rect 975 519 981 525
rect 987 519 993 525
rect 1011 519 1017 525
rect 1023 519 1029 525
rect 1035 519 1041 525
rect 1083 519 1089 525
rect 1095 519 1101 525
rect 1107 519 1113 525
rect 1131 519 1137 525
rect 1143 519 1149 525
rect 1155 519 1161 525
rect 1179 519 1185 525
rect 1191 519 1197 525
rect 1203 519 1209 525
rect 1227 519 1233 525
rect 1239 519 1245 525
rect 1251 519 1257 525
rect 1299 519 1305 525
rect 1311 519 1317 525
rect 1323 519 1329 525
rect 1347 519 1353 525
rect 1359 519 1365 525
rect 1371 519 1377 525
rect 1395 519 1401 525
rect 1407 519 1413 525
rect 1419 519 1425 525
rect 1443 519 1449 525
rect 1455 519 1461 525
rect 1467 519 1473 525
rect 3 423 9 429
rect 15 423 21 429
rect 27 423 33 429
rect 51 423 57 429
rect 63 423 69 429
rect 75 423 81 429
rect 99 423 105 429
rect 111 423 117 429
rect 123 423 129 429
rect 147 423 153 429
rect 159 423 165 429
rect 171 423 177 429
rect 219 423 225 429
rect 231 423 237 429
rect 243 423 249 429
rect 267 423 273 429
rect 279 423 285 429
rect 291 423 297 429
rect 315 423 321 429
rect 327 423 333 429
rect 339 423 345 429
rect 363 423 369 429
rect 375 423 381 429
rect 387 423 393 429
rect 435 423 441 429
rect 447 423 453 429
rect 459 423 465 429
rect 483 423 489 429
rect 495 423 501 429
rect 507 423 513 429
rect 531 423 537 429
rect 543 423 549 429
rect 555 423 561 429
rect 579 423 585 429
rect 591 423 597 429
rect 603 423 609 429
rect 651 423 657 429
rect 663 423 669 429
rect 675 423 681 429
rect 699 423 705 429
rect 711 423 717 429
rect 723 423 729 429
rect 747 423 753 429
rect 759 423 765 429
rect 771 423 777 429
rect 795 423 801 429
rect 807 423 813 429
rect 819 423 825 429
rect 867 423 873 429
rect 879 423 885 429
rect 891 423 897 429
rect 903 423 909 429
rect 915 423 921 429
rect 927 423 933 429
rect 939 423 945 429
rect 963 423 969 429
rect 975 423 981 429
rect 987 423 993 429
rect 1011 423 1017 429
rect 1023 423 1029 429
rect 1035 423 1041 429
rect 1083 423 1089 429
rect 1095 423 1101 429
rect 1107 423 1113 429
rect 1131 423 1137 429
rect 1143 423 1149 429
rect 1155 423 1161 429
rect 1179 423 1185 429
rect 1191 423 1197 429
rect 1203 423 1209 429
rect 1227 423 1233 429
rect 1239 423 1245 429
rect 1251 423 1257 429
rect 1299 423 1305 429
rect 1311 423 1317 429
rect 1323 423 1329 429
rect 1347 423 1353 429
rect 1359 423 1365 429
rect 1371 423 1377 429
rect 1395 423 1401 429
rect 1407 423 1413 429
rect 1419 423 1425 429
rect 1443 423 1449 429
rect 1455 423 1461 429
rect 1467 423 1473 429
rect 3 303 9 309
rect 15 303 21 309
rect 27 303 33 309
rect 51 303 57 309
rect 63 303 69 309
rect 75 303 81 309
rect 99 303 105 309
rect 111 303 117 309
rect 123 303 129 309
rect 147 303 153 309
rect 159 303 165 309
rect 171 303 177 309
rect 219 303 225 309
rect 231 303 237 309
rect 243 303 249 309
rect 267 303 273 309
rect 279 303 285 309
rect 291 303 297 309
rect 315 303 321 309
rect 327 303 333 309
rect 339 303 345 309
rect 363 303 369 309
rect 375 303 381 309
rect 387 303 393 309
rect 435 303 441 309
rect 447 303 453 309
rect 459 303 465 309
rect 483 303 489 309
rect 495 303 501 309
rect 507 303 513 309
rect 531 303 537 309
rect 543 303 549 309
rect 555 303 561 309
rect 579 303 585 309
rect 591 303 597 309
rect 603 303 609 309
rect 651 303 657 309
rect 663 303 669 309
rect 675 303 681 309
rect 699 303 705 309
rect 711 303 717 309
rect 723 303 729 309
rect 747 303 753 309
rect 759 303 765 309
rect 771 303 777 309
rect 795 303 801 309
rect 807 303 813 309
rect 819 303 825 309
rect 867 303 873 309
rect 915 303 921 309
rect 927 303 933 309
rect 939 303 945 309
rect 963 303 969 309
rect 975 303 981 309
rect 987 303 993 309
rect 1011 303 1017 309
rect 1023 303 1029 309
rect 1035 303 1041 309
rect 1083 303 1089 309
rect 1095 303 1101 309
rect 1107 303 1113 309
rect 1131 303 1137 309
rect 1143 303 1149 309
rect 1155 303 1161 309
rect 1179 303 1185 309
rect 1191 303 1197 309
rect 1203 303 1209 309
rect 1227 303 1233 309
rect 1239 303 1245 309
rect 1251 303 1257 309
rect 1299 303 1305 309
rect 1311 303 1317 309
rect 1323 303 1329 309
rect 1347 303 1353 309
rect 1359 303 1365 309
rect 1371 303 1377 309
rect 1395 303 1401 309
rect 1407 303 1413 309
rect 1419 303 1425 309
rect 1443 303 1449 309
rect 1455 303 1461 309
rect 1467 303 1473 309
rect 3 63 9 69
rect 15 63 21 69
rect 27 63 33 69
rect 51 63 57 69
rect 63 63 69 69
rect 75 63 81 69
rect 99 63 105 69
rect 111 63 117 69
rect 123 63 129 69
rect 147 63 153 69
rect 159 63 165 69
rect 171 63 177 69
rect 219 63 225 69
rect 231 63 237 69
rect 243 63 249 69
rect 267 63 273 69
rect 279 63 285 69
rect 291 63 297 69
rect 315 63 321 69
rect 327 63 333 69
rect 339 63 345 69
rect 363 63 369 69
rect 375 63 381 69
rect 387 63 393 69
rect 435 63 441 69
rect 447 63 453 69
rect 459 63 465 69
rect 483 63 489 69
rect 495 63 501 69
rect 507 63 513 69
rect 531 63 537 69
rect 543 63 549 69
rect 555 63 561 69
rect 579 63 585 69
rect 591 63 597 69
rect 603 63 609 69
rect 651 63 657 69
rect 663 63 669 69
rect 675 63 681 69
rect 699 63 705 69
rect 711 63 717 69
rect 723 63 729 69
rect 747 63 753 69
rect 759 63 765 69
rect 771 63 777 69
rect 795 63 801 69
rect 807 63 813 69
rect 819 63 825 69
rect 867 63 873 69
rect 879 63 885 69
rect 891 63 897 69
rect 915 63 921 69
rect 927 63 933 69
rect 939 63 945 69
rect 963 63 969 69
rect 975 63 981 69
rect 987 63 993 69
rect 1011 63 1017 69
rect 1023 63 1029 69
rect 1035 63 1041 69
rect 1083 63 1089 69
rect 1095 63 1101 69
rect 1107 63 1113 69
rect 1131 63 1137 69
rect 1143 63 1149 69
rect 1155 63 1161 69
rect 1179 63 1185 69
rect 1191 63 1197 69
rect 1203 63 1209 69
rect 1227 63 1233 69
rect 1239 63 1245 69
rect 1251 63 1257 69
rect 1299 63 1305 69
rect 1311 63 1317 69
rect 1323 63 1329 69
rect 1347 63 1353 69
rect 1359 63 1365 69
rect 1371 63 1377 69
rect 1395 63 1401 69
rect 1407 63 1413 69
rect 1419 63 1425 69
rect 1443 63 1449 69
rect 1455 63 1461 69
rect 1467 63 1473 69
<< metal1 >>
rect -60 621 1536 624
rect -60 615 -57 621
rect -51 615 -45 621
rect -39 615 -33 621
rect -27 615 -21 621
rect -15 615 -9 621
rect -3 615 3 621
rect 9 615 15 621
rect 21 615 27 621
rect 33 615 39 621
rect 45 615 51 621
rect 57 615 63 621
rect 69 615 75 621
rect 81 615 87 621
rect 93 615 99 621
rect 105 615 111 621
rect 117 615 123 621
rect 129 615 135 621
rect 141 615 147 621
rect 153 615 159 621
rect 165 615 171 621
rect 177 615 183 621
rect 189 615 195 621
rect 201 615 207 621
rect 213 615 219 621
rect 225 615 231 621
rect 237 615 243 621
rect 249 615 255 621
rect 261 615 267 621
rect 273 615 279 621
rect 285 615 291 621
rect 297 615 303 621
rect 309 615 315 621
rect 321 615 327 621
rect 333 615 339 621
rect 345 615 351 621
rect 357 615 363 621
rect 369 615 375 621
rect 381 615 387 621
rect 393 615 399 621
rect 405 615 411 621
rect 417 615 423 621
rect 429 615 435 621
rect 441 615 447 621
rect 453 615 459 621
rect 465 615 471 621
rect 477 615 483 621
rect 489 615 495 621
rect 501 615 507 621
rect 513 615 519 621
rect 525 615 531 621
rect 537 615 543 621
rect 549 615 555 621
rect 561 615 567 621
rect 573 615 579 621
rect 585 615 591 621
rect 597 615 603 621
rect 609 615 615 621
rect 621 615 627 621
rect 633 615 639 621
rect 645 615 651 621
rect 657 615 663 621
rect 669 615 675 621
rect 681 615 687 621
rect 693 615 699 621
rect 705 615 711 621
rect 717 615 723 621
rect 729 615 735 621
rect 741 615 747 621
rect 753 615 759 621
rect 765 615 771 621
rect 777 615 783 621
rect 789 615 795 621
rect 801 615 807 621
rect 813 615 819 621
rect 825 615 831 621
rect 837 615 843 621
rect 849 615 855 621
rect 861 615 867 621
rect 873 615 879 621
rect 885 615 891 621
rect 897 615 903 621
rect 909 615 915 621
rect 921 615 927 621
rect 933 615 939 621
rect 945 615 951 621
rect 957 615 963 621
rect 969 615 975 621
rect 981 615 987 621
rect 993 615 999 621
rect 1005 615 1011 621
rect 1017 615 1023 621
rect 1029 615 1035 621
rect 1041 615 1047 621
rect 1053 615 1059 621
rect 1065 615 1071 621
rect 1077 615 1083 621
rect 1089 615 1095 621
rect 1101 615 1107 621
rect 1113 615 1119 621
rect 1125 615 1131 621
rect 1137 615 1143 621
rect 1149 615 1155 621
rect 1161 615 1167 621
rect 1173 615 1179 621
rect 1185 615 1191 621
rect 1197 615 1203 621
rect 1209 615 1215 621
rect 1221 615 1227 621
rect 1233 615 1239 621
rect 1245 615 1251 621
rect 1257 615 1263 621
rect 1269 615 1275 621
rect 1281 615 1287 621
rect 1293 615 1299 621
rect 1305 615 1311 621
rect 1317 615 1323 621
rect 1329 615 1335 621
rect 1341 615 1347 621
rect 1353 615 1359 621
rect 1365 615 1371 621
rect 1377 615 1383 621
rect 1389 615 1395 621
rect 1401 615 1407 621
rect 1413 615 1419 621
rect 1425 615 1431 621
rect 1437 615 1443 621
rect 1449 615 1455 621
rect 1461 615 1467 621
rect 1473 615 1479 621
rect 1485 615 1491 621
rect 1497 615 1503 621
rect 1509 615 1515 621
rect 1521 615 1527 621
rect 1533 615 1536 621
rect -60 612 1536 615
rect -60 609 -48 612
rect -60 603 -57 609
rect -51 603 -48 609
rect -60 597 -48 603
rect 1524 609 1536 612
rect 1524 603 1527 609
rect 1533 603 1536 609
rect -60 591 -57 597
rect -51 591 -48 597
rect -60 585 -48 591
rect -60 579 -57 585
rect -51 579 -48 585
rect -60 573 -48 579
rect -60 567 -57 573
rect -51 567 -48 573
rect -60 561 -48 567
rect -60 555 -57 561
rect -51 555 -48 561
rect -60 549 -48 555
rect -60 543 -57 549
rect -51 543 -48 549
rect -60 537 -48 543
rect -60 531 -57 537
rect -51 531 -48 537
rect -60 525 -48 531
rect -60 519 -57 525
rect -51 519 -48 525
rect -60 513 -48 519
rect -60 507 -57 513
rect -51 507 -48 513
rect -60 501 -48 507
rect -60 495 -57 501
rect -51 495 -48 501
rect -60 489 -48 495
rect -60 483 -57 489
rect -51 483 -48 489
rect -60 477 -48 483
rect -60 471 -57 477
rect -51 471 -48 477
rect -60 465 -48 471
rect -60 459 -57 465
rect -51 459 -48 465
rect -60 453 -48 459
rect -60 447 -57 453
rect -51 447 -48 453
rect -60 441 -48 447
rect -60 435 -57 441
rect -51 435 -48 441
rect -60 429 -48 435
rect -60 423 -57 429
rect -51 423 -48 429
rect -60 417 -48 423
rect -60 411 -57 417
rect -51 411 -48 417
rect -60 405 -48 411
rect -60 399 -57 405
rect -51 399 -48 405
rect -60 393 -48 399
rect -60 387 -57 393
rect -51 387 -48 393
rect -60 381 -48 387
rect -60 375 -57 381
rect -51 375 -48 381
rect -60 369 -48 375
rect -60 363 -57 369
rect -51 363 -48 369
rect -60 357 -48 363
rect -60 351 -57 357
rect -51 351 -48 357
rect -60 345 -48 351
rect -36 597 1512 600
rect -36 591 -33 597
rect -27 591 -21 597
rect -15 591 -9 597
rect -3 591 3 597
rect 9 591 15 597
rect 21 591 27 597
rect 33 591 39 597
rect 45 591 51 597
rect 57 591 63 597
rect 69 591 75 597
rect 81 591 87 597
rect 93 591 99 597
rect 105 591 111 597
rect 117 591 123 597
rect 129 591 135 597
rect 141 591 147 597
rect 153 591 159 597
rect 165 591 171 597
rect 177 591 183 597
rect 189 591 195 597
rect 201 591 207 597
rect 213 591 219 597
rect 225 591 231 597
rect 237 591 243 597
rect 249 591 255 597
rect 261 591 267 597
rect 273 591 279 597
rect 285 591 291 597
rect 297 591 303 597
rect 309 591 315 597
rect 321 591 327 597
rect 333 591 339 597
rect 345 591 351 597
rect 357 591 363 597
rect 369 591 375 597
rect 381 591 387 597
rect 393 591 399 597
rect 405 591 411 597
rect 417 591 423 597
rect 429 591 435 597
rect 441 591 447 597
rect 453 591 459 597
rect 465 591 471 597
rect 477 591 483 597
rect 489 591 495 597
rect 501 591 507 597
rect 513 591 519 597
rect 525 591 531 597
rect 537 591 543 597
rect 549 591 555 597
rect 561 591 567 597
rect 573 591 579 597
rect 585 591 591 597
rect 597 591 603 597
rect 609 591 615 597
rect 621 591 627 597
rect 633 591 639 597
rect 645 591 651 597
rect 657 591 663 597
rect 669 591 675 597
rect 681 591 687 597
rect 693 591 699 597
rect 705 591 711 597
rect 717 591 723 597
rect 729 591 735 597
rect 741 591 747 597
rect 753 591 759 597
rect 765 591 771 597
rect 777 591 783 597
rect 789 591 795 597
rect 801 591 807 597
rect 813 591 819 597
rect 825 591 831 597
rect 837 591 843 597
rect 849 591 855 597
rect 861 591 867 597
rect 873 591 879 597
rect 885 591 891 597
rect 897 591 903 597
rect 909 591 915 597
rect 921 591 927 597
rect 933 591 939 597
rect 945 591 951 597
rect 957 591 963 597
rect 969 591 975 597
rect 981 591 987 597
rect 993 591 999 597
rect 1005 591 1011 597
rect 1017 591 1023 597
rect 1029 591 1035 597
rect 1041 591 1047 597
rect 1053 591 1059 597
rect 1065 591 1071 597
rect 1077 591 1083 597
rect 1089 591 1095 597
rect 1101 591 1107 597
rect 1113 591 1119 597
rect 1125 591 1131 597
rect 1137 591 1143 597
rect 1149 591 1155 597
rect 1161 591 1167 597
rect 1173 591 1179 597
rect 1185 591 1191 597
rect 1197 591 1203 597
rect 1209 591 1215 597
rect 1221 591 1227 597
rect 1233 591 1239 597
rect 1245 591 1251 597
rect 1257 591 1263 597
rect 1269 591 1275 597
rect 1281 591 1287 597
rect 1293 591 1299 597
rect 1305 591 1311 597
rect 1317 591 1323 597
rect 1329 591 1335 597
rect 1341 591 1347 597
rect 1353 591 1359 597
rect 1365 591 1371 597
rect 1377 591 1383 597
rect 1389 591 1395 597
rect 1401 591 1407 597
rect 1413 591 1419 597
rect 1425 591 1431 597
rect 1437 591 1443 597
rect 1449 591 1455 597
rect 1461 591 1467 597
rect 1473 591 1479 597
rect 1485 591 1491 597
rect 1497 591 1503 597
rect 1509 591 1512 597
rect -36 588 1512 591
rect -36 585 -24 588
rect -36 579 -33 585
rect -27 579 -24 585
rect -36 573 -24 579
rect -36 567 -33 573
rect -27 567 -24 573
rect -36 561 -24 567
rect -36 555 -33 561
rect -27 555 -24 561
rect -36 549 -24 555
rect -36 543 -33 549
rect -27 543 -24 549
rect -36 537 -24 543
rect -12 573 0 588
rect -12 567 -9 573
rect -3 567 0 573
rect -12 561 0 567
rect -12 555 -9 561
rect -3 555 0 561
rect -12 549 0 555
rect -12 543 -9 549
rect -3 543 0 549
rect -12 540 0 543
rect 12 573 24 576
rect 12 567 15 573
rect 21 567 24 573
rect 12 561 24 567
rect 12 555 15 561
rect 21 555 24 561
rect 12 549 24 555
rect 12 543 15 549
rect 21 543 24 549
rect 12 540 24 543
rect 36 573 48 588
rect 36 567 39 573
rect 45 567 48 573
rect 36 561 48 567
rect 36 555 39 561
rect 45 555 48 561
rect 36 549 48 555
rect 36 543 39 549
rect 45 543 48 549
rect 36 540 48 543
rect 60 573 72 576
rect 60 567 63 573
rect 69 567 72 573
rect 60 561 72 567
rect 60 555 63 561
rect 69 555 72 561
rect 60 549 72 555
rect 60 543 63 549
rect 69 543 72 549
rect 60 540 72 543
rect 84 573 96 588
rect 84 567 87 573
rect 93 567 96 573
rect 84 561 96 567
rect 84 555 87 561
rect 93 555 96 561
rect 84 549 96 555
rect 84 543 87 549
rect 93 543 96 549
rect 84 540 96 543
rect 108 573 120 576
rect 108 567 111 573
rect 117 567 120 573
rect 108 561 120 567
rect 108 555 111 561
rect 117 555 120 561
rect 108 549 120 555
rect 108 543 111 549
rect 117 543 120 549
rect 108 540 120 543
rect 132 573 144 588
rect 132 567 135 573
rect 141 567 144 573
rect 132 561 144 567
rect 132 555 135 561
rect 141 555 144 561
rect 132 549 144 555
rect 132 543 135 549
rect 141 543 144 549
rect 132 540 144 543
rect 156 573 168 576
rect 156 567 159 573
rect 165 567 168 573
rect 156 561 168 567
rect 156 555 159 561
rect 165 555 168 561
rect 156 549 168 555
rect 156 543 159 549
rect 165 543 168 549
rect 156 540 168 543
rect 180 573 192 588
rect 180 567 183 573
rect 189 567 192 573
rect 180 561 192 567
rect 180 555 183 561
rect 189 555 192 561
rect 180 549 192 555
rect 180 543 183 549
rect 189 543 192 549
rect 180 540 192 543
rect 204 573 216 588
rect 204 567 207 573
rect 213 567 216 573
rect 204 561 216 567
rect 204 555 207 561
rect 213 555 216 561
rect 204 549 216 555
rect 204 543 207 549
rect 213 543 216 549
rect 204 540 216 543
rect 252 573 264 576
rect 252 567 255 573
rect 261 567 264 573
rect 252 561 264 567
rect 252 555 255 561
rect 261 555 264 561
rect 252 549 264 555
rect 252 543 255 549
rect 261 543 264 549
rect 252 540 264 543
rect 300 573 312 588
rect 300 567 303 573
rect 309 567 312 573
rect 300 561 312 567
rect 300 555 303 561
rect 309 555 312 561
rect 300 549 312 555
rect 300 543 303 549
rect 309 543 312 549
rect 300 540 312 543
rect 348 573 360 576
rect 348 567 351 573
rect 357 567 360 573
rect 348 561 360 567
rect 348 555 351 561
rect 357 555 360 561
rect 348 549 360 555
rect 348 543 351 549
rect 357 543 360 549
rect 348 540 360 543
rect 396 573 408 588
rect 396 567 399 573
rect 405 567 408 573
rect 396 561 408 567
rect 396 555 399 561
rect 405 555 408 561
rect 396 549 408 555
rect 396 543 399 549
rect 405 543 408 549
rect 396 540 408 543
rect 420 573 432 588
rect 420 567 423 573
rect 429 567 432 573
rect 420 561 432 567
rect 420 555 423 561
rect 429 555 432 561
rect 420 549 432 555
rect 420 543 423 549
rect 429 543 432 549
rect 420 540 432 543
rect 468 573 480 576
rect 468 567 471 573
rect 477 567 480 573
rect 468 561 480 567
rect 468 555 471 561
rect 477 555 480 561
rect 468 549 480 555
rect 468 543 471 549
rect 477 543 480 549
rect 468 540 480 543
rect 516 573 528 588
rect 516 567 519 573
rect 525 567 528 573
rect 516 561 528 567
rect 516 555 519 561
rect 525 555 528 561
rect 516 549 528 555
rect 516 543 519 549
rect 525 543 528 549
rect 516 540 528 543
rect 564 573 576 576
rect 564 567 567 573
rect 573 567 576 573
rect 564 561 576 567
rect 564 555 567 561
rect 573 555 576 561
rect 564 549 576 555
rect 564 543 567 549
rect 573 543 576 549
rect 564 540 576 543
rect 612 573 624 588
rect 612 567 615 573
rect 621 567 624 573
rect 612 561 624 567
rect 612 555 615 561
rect 621 555 624 561
rect 612 549 624 555
rect 612 543 615 549
rect 621 543 624 549
rect 612 540 624 543
rect 636 573 648 588
rect 636 567 639 573
rect 645 567 648 573
rect 636 561 648 567
rect 636 555 639 561
rect 645 555 648 561
rect 636 549 648 555
rect 636 543 639 549
rect 645 543 648 549
rect 636 540 648 543
rect 828 573 840 576
rect 828 567 831 573
rect 837 567 840 573
rect 828 561 840 567
rect 828 555 831 561
rect 837 555 840 561
rect 828 549 840 555
rect 828 543 831 549
rect 837 543 840 549
rect 828 540 840 543
rect 852 573 864 588
rect 852 567 855 573
rect 861 567 864 573
rect 852 561 864 567
rect 852 555 855 561
rect 861 555 864 561
rect 852 549 864 555
rect 852 543 855 549
rect 861 543 864 549
rect 852 540 864 543
rect 1044 573 1056 576
rect 1044 567 1047 573
rect 1053 567 1056 573
rect 1044 561 1056 567
rect 1044 555 1047 561
rect 1053 555 1056 561
rect 1044 549 1056 555
rect 1044 543 1047 549
rect 1053 543 1056 549
rect 1044 540 1056 543
rect 1068 573 1080 588
rect 1068 567 1071 573
rect 1077 567 1080 573
rect 1068 561 1080 567
rect 1068 555 1071 561
rect 1077 555 1080 561
rect 1068 549 1080 555
rect 1068 543 1071 549
rect 1077 543 1080 549
rect 1068 540 1080 543
rect 1092 573 1104 576
rect 1092 567 1095 573
rect 1101 567 1104 573
rect 1092 561 1104 567
rect 1092 555 1095 561
rect 1101 555 1104 561
rect 1092 549 1104 555
rect 1092 543 1095 549
rect 1101 543 1104 549
rect 1092 540 1104 543
rect 1116 573 1128 588
rect 1116 567 1119 573
rect 1125 567 1128 573
rect 1116 561 1128 567
rect 1116 555 1119 561
rect 1125 555 1128 561
rect 1116 549 1128 555
rect 1116 543 1119 549
rect 1125 543 1128 549
rect 1116 540 1128 543
rect 1140 573 1152 576
rect 1140 567 1143 573
rect 1149 567 1152 573
rect 1140 561 1152 567
rect 1140 555 1143 561
rect 1149 555 1152 561
rect 1140 549 1152 555
rect 1140 543 1143 549
rect 1149 543 1152 549
rect 1140 540 1152 543
rect 1164 573 1176 588
rect 1164 567 1167 573
rect 1173 567 1176 573
rect 1164 561 1176 567
rect 1164 555 1167 561
rect 1173 555 1176 561
rect 1164 549 1176 555
rect 1164 543 1167 549
rect 1173 543 1176 549
rect 1164 540 1176 543
rect 1188 573 1200 576
rect 1188 567 1191 573
rect 1197 567 1200 573
rect 1188 561 1200 567
rect 1188 555 1191 561
rect 1197 555 1200 561
rect 1188 549 1200 555
rect 1188 543 1191 549
rect 1197 543 1200 549
rect 1188 540 1200 543
rect 1212 573 1224 588
rect 1212 567 1215 573
rect 1221 567 1224 573
rect 1212 561 1224 567
rect 1212 555 1215 561
rect 1221 555 1224 561
rect 1212 549 1224 555
rect 1212 543 1215 549
rect 1221 543 1224 549
rect 1212 540 1224 543
rect 1236 573 1248 576
rect 1236 567 1239 573
rect 1245 567 1248 573
rect 1236 561 1248 567
rect 1236 555 1239 561
rect 1245 555 1248 561
rect 1236 549 1248 555
rect 1236 543 1239 549
rect 1245 543 1248 549
rect 1236 540 1248 543
rect 1260 573 1272 588
rect 1260 567 1263 573
rect 1269 567 1272 573
rect 1260 561 1272 567
rect 1260 555 1263 561
rect 1269 555 1272 561
rect 1260 549 1272 555
rect 1260 543 1263 549
rect 1269 543 1272 549
rect 1260 540 1272 543
rect 1284 573 1296 588
rect 1284 567 1287 573
rect 1293 567 1296 573
rect 1284 561 1296 567
rect 1284 555 1287 561
rect 1293 555 1296 561
rect 1284 549 1296 555
rect 1284 543 1287 549
rect 1293 543 1296 549
rect 1284 540 1296 543
rect 1308 573 1320 576
rect 1308 567 1311 573
rect 1317 567 1320 573
rect 1308 561 1320 567
rect 1308 555 1311 561
rect 1317 555 1320 561
rect 1308 549 1320 555
rect 1308 543 1311 549
rect 1317 543 1320 549
rect 1308 540 1320 543
rect 1332 573 1344 588
rect 1332 567 1335 573
rect 1341 567 1344 573
rect 1332 561 1344 567
rect 1332 555 1335 561
rect 1341 555 1344 561
rect 1332 549 1344 555
rect 1332 543 1335 549
rect 1341 543 1344 549
rect 1332 540 1344 543
rect 1356 573 1368 576
rect 1356 567 1359 573
rect 1365 567 1368 573
rect 1356 561 1368 567
rect 1356 555 1359 561
rect 1365 555 1368 561
rect 1356 549 1368 555
rect 1356 543 1359 549
rect 1365 543 1368 549
rect 1356 540 1368 543
rect 1380 573 1392 588
rect 1380 567 1383 573
rect 1389 567 1392 573
rect 1380 561 1392 567
rect 1380 555 1383 561
rect 1389 555 1392 561
rect 1380 549 1392 555
rect 1380 543 1383 549
rect 1389 543 1392 549
rect 1380 540 1392 543
rect 1404 573 1416 576
rect 1404 567 1407 573
rect 1413 567 1416 573
rect 1404 561 1416 567
rect 1404 555 1407 561
rect 1413 555 1416 561
rect 1404 549 1416 555
rect 1404 543 1407 549
rect 1413 543 1416 549
rect 1404 540 1416 543
rect 1428 573 1440 588
rect 1428 567 1431 573
rect 1437 567 1440 573
rect 1428 561 1440 567
rect 1428 555 1431 561
rect 1437 555 1440 561
rect 1428 549 1440 555
rect 1428 543 1431 549
rect 1437 543 1440 549
rect 1428 540 1440 543
rect 1452 573 1464 576
rect 1452 567 1455 573
rect 1461 567 1464 573
rect 1452 561 1464 567
rect 1452 555 1455 561
rect 1461 555 1464 561
rect 1452 549 1464 555
rect 1452 543 1455 549
rect 1461 543 1464 549
rect 1452 540 1464 543
rect 1476 573 1488 588
rect 1476 567 1479 573
rect 1485 567 1488 573
rect 1476 561 1488 567
rect 1476 555 1479 561
rect 1485 555 1488 561
rect 1476 549 1488 555
rect 1476 543 1479 549
rect 1485 543 1488 549
rect 1476 540 1488 543
rect 1500 585 1512 588
rect 1500 579 1503 585
rect 1509 579 1512 585
rect 1500 573 1512 579
rect 1500 567 1503 573
rect 1509 567 1512 573
rect 1500 561 1512 567
rect 1500 555 1503 561
rect 1509 555 1512 561
rect 1500 549 1512 555
rect 1500 543 1503 549
rect 1509 543 1512 549
rect -36 531 -33 537
rect -27 531 -24 537
rect -36 525 -24 531
rect 1500 537 1512 543
rect 1500 531 1503 537
rect 1509 531 1512 537
rect -36 519 -33 525
rect -27 519 -24 525
rect -36 513 -24 519
rect 0 525 180 528
rect 0 519 3 525
rect 9 519 15 525
rect 21 519 27 525
rect 33 519 39 525
rect 45 519 51 525
rect 57 519 63 525
rect 69 519 75 525
rect 81 519 87 525
rect 93 519 99 525
rect 105 519 111 525
rect 117 519 123 525
rect 129 519 135 525
rect 141 519 147 525
rect 153 519 159 525
rect 165 519 171 525
rect 177 519 180 525
rect 0 516 180 519
rect 216 525 252 528
rect 216 519 219 525
rect 225 519 231 525
rect 237 519 243 525
rect 249 519 252 525
rect 216 516 252 519
rect 264 525 300 528
rect 264 519 267 525
rect 273 519 279 525
rect 285 519 291 525
rect 297 519 300 525
rect 264 516 300 519
rect 312 525 348 528
rect 312 519 315 525
rect 321 519 327 525
rect 333 519 339 525
rect 345 519 348 525
rect 312 516 348 519
rect 360 525 396 528
rect 360 519 363 525
rect 369 519 375 525
rect 381 519 387 525
rect 393 519 396 525
rect 360 516 396 519
rect 432 525 612 528
rect 432 519 435 525
rect 441 519 447 525
rect 453 519 459 525
rect 465 519 483 525
rect 489 519 495 525
rect 501 519 507 525
rect 513 519 519 525
rect 525 519 531 525
rect 537 519 543 525
rect 549 519 555 525
rect 561 519 579 525
rect 585 519 591 525
rect 597 519 603 525
rect 609 519 612 525
rect 432 516 612 519
rect 636 525 828 528
rect 636 519 639 525
rect 645 519 651 525
rect 657 519 663 525
rect 669 519 675 525
rect 681 519 699 525
rect 705 519 711 525
rect 717 519 723 525
rect 729 519 747 525
rect 753 519 759 525
rect 765 519 771 525
rect 777 519 795 525
rect 801 519 807 525
rect 813 519 819 525
rect 825 519 828 525
rect 636 516 828 519
rect 864 525 1044 528
rect 864 519 867 525
rect 873 519 879 525
rect 885 519 891 525
rect 897 519 903 525
rect 909 519 915 525
rect 921 519 927 525
rect 933 519 939 525
rect 945 519 963 525
rect 969 519 975 525
rect 981 519 987 525
rect 993 519 1011 525
rect 1017 519 1023 525
rect 1029 519 1035 525
rect 1041 519 1044 525
rect 864 516 1044 519
rect 1080 525 1260 528
rect 1080 519 1083 525
rect 1089 519 1095 525
rect 1101 519 1107 525
rect 1113 519 1119 525
rect 1125 519 1131 525
rect 1137 519 1143 525
rect 1149 519 1155 525
rect 1161 519 1167 525
rect 1173 519 1179 525
rect 1185 519 1191 525
rect 1197 519 1203 525
rect 1209 519 1215 525
rect 1221 519 1227 525
rect 1233 519 1239 525
rect 1245 519 1251 525
rect 1257 519 1260 525
rect 1080 516 1260 519
rect 1296 525 1476 528
rect 1296 519 1299 525
rect 1305 519 1311 525
rect 1317 519 1323 525
rect 1329 519 1335 525
rect 1341 519 1347 525
rect 1353 519 1359 525
rect 1365 519 1371 525
rect 1377 519 1383 525
rect 1389 519 1395 525
rect 1401 519 1407 525
rect 1413 519 1419 525
rect 1425 519 1431 525
rect 1437 519 1443 525
rect 1449 519 1455 525
rect 1461 519 1467 525
rect 1473 519 1476 525
rect 1296 516 1476 519
rect 1500 525 1512 531
rect 1500 519 1503 525
rect 1509 519 1512 525
rect -36 507 -33 513
rect -27 507 -24 513
rect -36 504 -24 507
rect 1500 513 1512 519
rect 1500 507 1503 513
rect 1509 507 1512 513
rect 1500 504 1512 507
rect -36 501 1512 504
rect -36 495 -33 501
rect -27 495 -21 501
rect -15 495 -9 501
rect -3 495 3 501
rect 9 495 15 501
rect 21 495 27 501
rect 33 495 39 501
rect 45 495 51 501
rect 57 495 63 501
rect 69 495 75 501
rect 81 495 87 501
rect 93 495 99 501
rect 105 495 111 501
rect 117 495 123 501
rect 129 495 135 501
rect 141 495 147 501
rect 153 495 159 501
rect 165 495 171 501
rect 177 495 183 501
rect 189 495 195 501
rect 201 495 207 501
rect 213 495 219 501
rect 225 495 231 501
rect 237 495 243 501
rect 249 495 255 501
rect 261 495 267 501
rect 273 495 279 501
rect 285 495 291 501
rect 297 495 303 501
rect 309 495 315 501
rect 321 495 327 501
rect 333 495 339 501
rect 345 495 351 501
rect 357 495 363 501
rect 369 495 375 501
rect 381 495 387 501
rect 393 495 399 501
rect 405 495 411 501
rect 417 495 423 501
rect 429 495 435 501
rect 441 495 447 501
rect 453 495 459 501
rect 465 495 471 501
rect 477 495 483 501
rect 489 495 495 501
rect 501 495 507 501
rect 513 495 519 501
rect 525 495 531 501
rect 537 495 543 501
rect 549 495 555 501
rect 561 495 567 501
rect 573 495 579 501
rect 585 495 591 501
rect 597 495 603 501
rect 609 495 615 501
rect 621 495 627 501
rect 633 495 639 501
rect 645 495 651 501
rect 657 495 663 501
rect 669 495 675 501
rect 681 495 687 501
rect 693 495 699 501
rect 705 495 711 501
rect 717 495 723 501
rect 729 495 735 501
rect 741 495 747 501
rect 753 495 759 501
rect 765 495 771 501
rect 777 495 783 501
rect 789 495 795 501
rect 801 495 807 501
rect 813 495 819 501
rect 825 495 831 501
rect 837 495 843 501
rect 849 495 855 501
rect 861 495 867 501
rect 873 495 879 501
rect 885 495 891 501
rect 897 495 903 501
rect 909 495 915 501
rect 921 495 927 501
rect 933 495 939 501
rect 945 495 951 501
rect 957 495 963 501
rect 969 495 975 501
rect 981 495 987 501
rect 993 495 999 501
rect 1005 495 1011 501
rect 1017 495 1023 501
rect 1029 495 1035 501
rect 1041 495 1047 501
rect 1053 495 1059 501
rect 1065 495 1071 501
rect 1077 495 1083 501
rect 1089 495 1095 501
rect 1101 495 1107 501
rect 1113 495 1119 501
rect 1125 495 1131 501
rect 1137 495 1143 501
rect 1149 495 1155 501
rect 1161 495 1167 501
rect 1173 495 1179 501
rect 1185 495 1191 501
rect 1197 495 1203 501
rect 1209 495 1215 501
rect 1221 495 1227 501
rect 1233 495 1239 501
rect 1245 495 1251 501
rect 1257 495 1263 501
rect 1269 495 1275 501
rect 1281 495 1287 501
rect 1293 495 1299 501
rect 1305 495 1311 501
rect 1317 495 1323 501
rect 1329 495 1335 501
rect 1341 495 1347 501
rect 1353 495 1359 501
rect 1365 495 1371 501
rect 1377 495 1383 501
rect 1389 495 1395 501
rect 1401 495 1407 501
rect 1413 495 1419 501
rect 1425 495 1431 501
rect 1437 495 1443 501
rect 1449 495 1455 501
rect 1461 495 1467 501
rect 1473 495 1479 501
rect 1485 495 1491 501
rect 1497 495 1503 501
rect 1509 495 1512 501
rect -36 492 1512 495
rect -36 489 -24 492
rect -36 483 -33 489
rect -27 483 -24 489
rect -36 477 -24 483
rect 1500 489 1512 492
rect 1500 483 1503 489
rect 1509 483 1512 489
rect -36 471 -33 477
rect -27 471 -24 477
rect -36 465 -24 471
rect -36 459 -33 465
rect -27 459 -24 465
rect -36 453 -24 459
rect -36 447 -33 453
rect -27 447 -24 453
rect -36 441 -24 447
rect -12 477 0 480
rect -12 471 -9 477
rect -3 471 0 477
rect -12 465 0 471
rect -12 459 -9 465
rect -3 459 0 465
rect -12 453 0 459
rect -12 447 -9 453
rect -3 447 0 453
rect -12 444 0 447
rect 12 477 24 480
rect 12 471 15 477
rect 21 471 24 477
rect 12 465 24 471
rect 12 459 15 465
rect 21 459 24 465
rect 12 453 24 459
rect 12 447 15 453
rect 21 447 24 453
rect 12 444 24 447
rect 36 477 48 480
rect 36 471 39 477
rect 45 471 48 477
rect 36 465 48 471
rect 36 459 39 465
rect 45 459 48 465
rect 36 453 48 459
rect 36 447 39 453
rect 45 447 48 453
rect 36 444 48 447
rect 60 477 72 480
rect 60 471 63 477
rect 69 471 72 477
rect 60 465 72 471
rect 60 459 63 465
rect 69 459 72 465
rect 60 453 72 459
rect 60 447 63 453
rect 69 447 72 453
rect 60 444 72 447
rect 84 477 96 480
rect 84 471 87 477
rect 93 471 96 477
rect 84 465 96 471
rect 84 459 87 465
rect 93 459 96 465
rect 84 453 96 459
rect 84 447 87 453
rect 93 447 96 453
rect 84 444 96 447
rect 108 477 120 480
rect 108 471 111 477
rect 117 471 120 477
rect 108 465 120 471
rect 108 459 111 465
rect 117 459 120 465
rect 108 453 120 459
rect 108 447 111 453
rect 117 447 120 453
rect 108 444 120 447
rect 132 477 144 480
rect 132 471 135 477
rect 141 471 144 477
rect 132 465 144 471
rect 132 459 135 465
rect 141 459 144 465
rect 132 453 144 459
rect 132 447 135 453
rect 141 447 144 453
rect 132 444 144 447
rect 156 477 168 480
rect 156 471 159 477
rect 165 471 168 477
rect 156 465 168 471
rect 156 459 159 465
rect 165 459 168 465
rect 156 453 168 459
rect 156 447 159 453
rect 165 447 168 453
rect 156 444 168 447
rect 180 477 192 480
rect 180 471 183 477
rect 189 471 192 477
rect 180 465 192 471
rect 180 459 183 465
rect 189 459 192 465
rect 180 453 192 459
rect 180 447 183 453
rect 189 447 192 453
rect 180 444 192 447
rect 204 477 216 480
rect 204 471 207 477
rect 213 471 216 477
rect 204 465 216 471
rect 204 459 207 465
rect 213 459 216 465
rect 204 453 216 459
rect 204 447 207 453
rect 213 447 216 453
rect 204 444 216 447
rect 252 477 264 480
rect 252 471 255 477
rect 261 471 264 477
rect 252 465 264 471
rect 252 459 255 465
rect 261 459 264 465
rect 252 453 264 459
rect 252 447 255 453
rect 261 447 264 453
rect 252 444 264 447
rect 300 477 312 480
rect 300 471 303 477
rect 309 471 312 477
rect 300 465 312 471
rect 300 459 303 465
rect 309 459 312 465
rect 300 453 312 459
rect 300 447 303 453
rect 309 447 312 453
rect 300 444 312 447
rect 348 477 360 480
rect 348 471 351 477
rect 357 471 360 477
rect 348 465 360 471
rect 348 459 351 465
rect 357 459 360 465
rect 348 453 360 459
rect 348 447 351 453
rect 357 447 360 453
rect 348 444 360 447
rect 396 477 408 480
rect 396 471 399 477
rect 405 471 408 477
rect 396 465 408 471
rect 396 459 399 465
rect 405 459 408 465
rect 396 453 408 459
rect 396 447 399 453
rect 405 447 408 453
rect 396 444 408 447
rect 420 477 432 480
rect 420 471 423 477
rect 429 471 432 477
rect 420 465 432 471
rect 420 459 423 465
rect 429 459 432 465
rect 420 453 432 459
rect 420 447 423 453
rect 429 447 432 453
rect 420 444 432 447
rect 468 477 480 480
rect 468 471 471 477
rect 477 471 480 477
rect 468 465 480 471
rect 468 459 471 465
rect 477 459 480 465
rect 468 453 480 459
rect 468 447 471 453
rect 477 447 480 453
rect 468 444 480 447
rect 516 477 528 480
rect 516 471 519 477
rect 525 471 528 477
rect 516 465 528 471
rect 516 459 519 465
rect 525 459 528 465
rect 516 453 528 459
rect 516 447 519 453
rect 525 447 528 453
rect 516 444 528 447
rect 564 477 576 480
rect 564 471 567 477
rect 573 471 576 477
rect 564 465 576 471
rect 564 459 567 465
rect 573 459 576 465
rect 564 453 576 459
rect 564 447 567 453
rect 573 447 576 453
rect 564 444 576 447
rect 612 477 624 480
rect 612 471 615 477
rect 621 471 624 477
rect 612 465 624 471
rect 612 459 615 465
rect 621 459 624 465
rect 612 453 624 459
rect 612 447 615 453
rect 621 447 624 453
rect 612 444 624 447
rect 636 477 648 480
rect 636 471 639 477
rect 645 471 648 477
rect 636 465 648 471
rect 636 459 639 465
rect 645 459 648 465
rect 636 453 648 459
rect 636 447 639 453
rect 645 447 648 453
rect 636 444 648 447
rect 828 477 840 480
rect 828 471 831 477
rect 837 471 840 477
rect 828 465 840 471
rect 828 459 831 465
rect 837 459 840 465
rect 828 453 840 459
rect 828 447 831 453
rect 837 447 840 453
rect 828 444 840 447
rect 852 477 864 480
rect 852 471 855 477
rect 861 471 864 477
rect 852 465 864 471
rect 852 459 855 465
rect 861 459 864 465
rect 852 453 864 459
rect 852 447 855 453
rect 861 447 864 453
rect 852 444 864 447
rect 1044 477 1056 480
rect 1044 471 1047 477
rect 1053 471 1056 477
rect 1044 465 1056 471
rect 1044 459 1047 465
rect 1053 459 1056 465
rect 1044 453 1056 459
rect 1044 447 1047 453
rect 1053 447 1056 453
rect 1044 444 1056 447
rect 1068 477 1080 480
rect 1068 471 1071 477
rect 1077 471 1080 477
rect 1068 465 1080 471
rect 1068 459 1071 465
rect 1077 459 1080 465
rect 1068 453 1080 459
rect 1068 447 1071 453
rect 1077 447 1080 453
rect 1068 444 1080 447
rect 1092 477 1104 480
rect 1092 471 1095 477
rect 1101 471 1104 477
rect 1092 465 1104 471
rect 1092 459 1095 465
rect 1101 459 1104 465
rect 1092 453 1104 459
rect 1092 447 1095 453
rect 1101 447 1104 453
rect 1092 444 1104 447
rect 1116 477 1128 480
rect 1116 471 1119 477
rect 1125 471 1128 477
rect 1116 465 1128 471
rect 1116 459 1119 465
rect 1125 459 1128 465
rect 1116 453 1128 459
rect 1116 447 1119 453
rect 1125 447 1128 453
rect 1116 444 1128 447
rect 1140 477 1152 480
rect 1140 471 1143 477
rect 1149 471 1152 477
rect 1140 465 1152 471
rect 1140 459 1143 465
rect 1149 459 1152 465
rect 1140 453 1152 459
rect 1140 447 1143 453
rect 1149 447 1152 453
rect 1140 444 1152 447
rect 1164 477 1176 480
rect 1164 471 1167 477
rect 1173 471 1176 477
rect 1164 465 1176 471
rect 1164 459 1167 465
rect 1173 459 1176 465
rect 1164 453 1176 459
rect 1164 447 1167 453
rect 1173 447 1176 453
rect 1164 444 1176 447
rect 1188 477 1200 480
rect 1188 471 1191 477
rect 1197 471 1200 477
rect 1188 465 1200 471
rect 1188 459 1191 465
rect 1197 459 1200 465
rect 1188 453 1200 459
rect 1188 447 1191 453
rect 1197 447 1200 453
rect 1188 444 1200 447
rect 1212 477 1224 480
rect 1212 471 1215 477
rect 1221 471 1224 477
rect 1212 465 1224 471
rect 1212 459 1215 465
rect 1221 459 1224 465
rect 1212 453 1224 459
rect 1212 447 1215 453
rect 1221 447 1224 453
rect 1212 444 1224 447
rect 1236 477 1248 480
rect 1236 471 1239 477
rect 1245 471 1248 477
rect 1236 465 1248 471
rect 1236 459 1239 465
rect 1245 459 1248 465
rect 1236 453 1248 459
rect 1236 447 1239 453
rect 1245 447 1248 453
rect 1236 444 1248 447
rect 1260 477 1272 480
rect 1260 471 1263 477
rect 1269 471 1272 477
rect 1260 465 1272 471
rect 1260 459 1263 465
rect 1269 459 1272 465
rect 1260 453 1272 459
rect 1260 447 1263 453
rect 1269 447 1272 453
rect 1260 444 1272 447
rect 1284 477 1296 480
rect 1284 471 1287 477
rect 1293 471 1296 477
rect 1284 465 1296 471
rect 1284 459 1287 465
rect 1293 459 1296 465
rect 1284 453 1296 459
rect 1284 447 1287 453
rect 1293 447 1296 453
rect 1284 444 1296 447
rect 1308 477 1320 480
rect 1308 471 1311 477
rect 1317 471 1320 477
rect 1308 465 1320 471
rect 1308 459 1311 465
rect 1317 459 1320 465
rect 1308 453 1320 459
rect 1308 447 1311 453
rect 1317 447 1320 453
rect 1308 444 1320 447
rect 1332 477 1344 480
rect 1332 471 1335 477
rect 1341 471 1344 477
rect 1332 465 1344 471
rect 1332 459 1335 465
rect 1341 459 1344 465
rect 1332 453 1344 459
rect 1332 447 1335 453
rect 1341 447 1344 453
rect 1332 444 1344 447
rect 1356 477 1368 480
rect 1356 471 1359 477
rect 1365 471 1368 477
rect 1356 465 1368 471
rect 1356 459 1359 465
rect 1365 459 1368 465
rect 1356 453 1368 459
rect 1356 447 1359 453
rect 1365 447 1368 453
rect 1356 444 1368 447
rect 1380 477 1392 480
rect 1380 471 1383 477
rect 1389 471 1392 477
rect 1380 465 1392 471
rect 1380 459 1383 465
rect 1389 459 1392 465
rect 1380 453 1392 459
rect 1380 447 1383 453
rect 1389 447 1392 453
rect 1380 444 1392 447
rect 1404 477 1416 480
rect 1404 471 1407 477
rect 1413 471 1416 477
rect 1404 465 1416 471
rect 1404 459 1407 465
rect 1413 459 1416 465
rect 1404 453 1416 459
rect 1404 447 1407 453
rect 1413 447 1416 453
rect 1404 444 1416 447
rect 1428 477 1440 480
rect 1428 471 1431 477
rect 1437 471 1440 477
rect 1428 465 1440 471
rect 1428 459 1431 465
rect 1437 459 1440 465
rect 1428 453 1440 459
rect 1428 447 1431 453
rect 1437 447 1440 453
rect 1428 444 1440 447
rect 1452 477 1464 480
rect 1452 471 1455 477
rect 1461 471 1464 477
rect 1452 465 1464 471
rect 1452 459 1455 465
rect 1461 459 1464 465
rect 1452 453 1464 459
rect 1452 447 1455 453
rect 1461 447 1464 453
rect 1452 444 1464 447
rect 1476 477 1488 480
rect 1476 471 1479 477
rect 1485 471 1488 477
rect 1476 465 1488 471
rect 1476 459 1479 465
rect 1485 459 1488 465
rect 1476 453 1488 459
rect 1476 447 1479 453
rect 1485 447 1488 453
rect 1476 444 1488 447
rect 1500 477 1512 483
rect 1500 471 1503 477
rect 1509 471 1512 477
rect 1500 465 1512 471
rect 1500 459 1503 465
rect 1509 459 1512 465
rect 1500 453 1512 459
rect 1500 447 1503 453
rect 1509 447 1512 453
rect -36 435 -33 441
rect -27 435 -24 441
rect -36 429 -24 435
rect 1500 441 1512 447
rect 1500 435 1503 441
rect 1509 435 1512 441
rect -36 423 -33 429
rect -27 423 -24 429
rect -36 417 -24 423
rect 0 429 36 432
rect 0 423 3 429
rect 9 423 15 429
rect 21 423 27 429
rect 33 423 36 429
rect 0 420 36 423
rect 48 429 84 432
rect 48 423 51 429
rect 57 423 63 429
rect 69 423 75 429
rect 81 423 84 429
rect 48 420 84 423
rect 96 429 132 432
rect 96 423 99 429
rect 105 423 111 429
rect 117 423 123 429
rect 129 423 132 429
rect 96 420 132 423
rect 144 429 180 432
rect 144 423 147 429
rect 153 423 159 429
rect 165 423 171 429
rect 177 423 180 429
rect 144 420 180 423
rect 216 429 252 432
rect 216 423 219 429
rect 225 423 231 429
rect 237 423 243 429
rect 249 423 252 429
rect 216 420 252 423
rect 264 429 300 432
rect 264 423 267 429
rect 273 423 279 429
rect 285 423 291 429
rect 297 423 300 429
rect 264 420 300 423
rect 312 429 348 432
rect 312 423 315 429
rect 321 423 327 429
rect 333 423 339 429
rect 345 423 348 429
rect 312 420 348 423
rect 360 429 396 432
rect 360 423 363 429
rect 369 423 375 429
rect 381 423 387 429
rect 393 423 396 429
rect 360 420 396 423
rect 432 429 468 432
rect 432 423 435 429
rect 441 423 447 429
rect 453 423 459 429
rect 465 423 468 429
rect 432 420 468 423
rect 480 429 516 432
rect 480 423 483 429
rect 489 423 495 429
rect 501 423 507 429
rect 513 423 516 429
rect 480 420 516 423
rect 528 429 564 432
rect 528 423 531 429
rect 537 423 543 429
rect 549 423 555 429
rect 561 423 564 429
rect 528 420 564 423
rect 576 429 612 432
rect 576 423 579 429
rect 585 423 591 429
rect 597 423 603 429
rect 609 423 612 429
rect 576 420 612 423
rect 636 429 684 432
rect 636 423 639 429
rect 645 423 651 429
rect 657 423 663 429
rect 669 423 675 429
rect 681 423 684 429
rect 636 420 684 423
rect 696 429 732 432
rect 696 423 699 429
rect 705 423 711 429
rect 717 423 723 429
rect 729 423 732 429
rect 696 420 732 423
rect 744 429 780 432
rect 744 423 747 429
rect 753 423 759 429
rect 765 423 771 429
rect 777 423 780 429
rect 744 420 780 423
rect 792 429 840 432
rect 792 423 795 429
rect 801 423 807 429
rect 813 423 819 429
rect 825 423 831 429
rect 837 423 840 429
rect 792 420 840 423
rect 864 429 1044 432
rect 864 423 867 429
rect 873 423 879 429
rect 885 423 891 429
rect 897 423 903 429
rect 909 423 915 429
rect 921 423 927 429
rect 933 423 939 429
rect 945 423 963 429
rect 969 423 975 429
rect 981 423 987 429
rect 993 423 1011 429
rect 1017 423 1023 429
rect 1029 423 1035 429
rect 1041 423 1044 429
rect 864 420 1044 423
rect 1080 429 1116 432
rect 1080 423 1083 429
rect 1089 423 1095 429
rect 1101 423 1107 429
rect 1113 423 1116 429
rect 1080 420 1116 423
rect 1128 429 1164 432
rect 1128 423 1131 429
rect 1137 423 1143 429
rect 1149 423 1155 429
rect 1161 423 1164 429
rect 1128 420 1164 423
rect 1176 429 1212 432
rect 1176 423 1179 429
rect 1185 423 1191 429
rect 1197 423 1203 429
rect 1209 423 1212 429
rect 1176 420 1212 423
rect 1224 429 1260 432
rect 1224 423 1227 429
rect 1233 423 1239 429
rect 1245 423 1251 429
rect 1257 423 1260 429
rect 1224 420 1260 423
rect 1296 429 1332 432
rect 1296 423 1299 429
rect 1305 423 1311 429
rect 1317 423 1323 429
rect 1329 423 1332 429
rect 1296 420 1332 423
rect 1344 429 1380 432
rect 1344 423 1347 429
rect 1353 423 1359 429
rect 1365 423 1371 429
rect 1377 423 1380 429
rect 1344 420 1380 423
rect 1392 429 1428 432
rect 1392 423 1395 429
rect 1401 423 1407 429
rect 1413 423 1419 429
rect 1425 423 1428 429
rect 1392 420 1428 423
rect 1440 429 1476 432
rect 1440 423 1443 429
rect 1449 423 1455 429
rect 1461 423 1467 429
rect 1473 423 1476 429
rect 1440 420 1476 423
rect 1500 429 1512 435
rect 1500 423 1503 429
rect 1509 423 1512 429
rect -36 411 -33 417
rect -27 411 -24 417
rect -36 408 -24 411
rect 1500 417 1512 423
rect 1500 411 1503 417
rect 1509 411 1512 417
rect 1500 408 1512 411
rect -36 405 1512 408
rect -36 399 -33 405
rect -27 399 -21 405
rect -15 399 -9 405
rect -3 399 3 405
rect 9 399 15 405
rect 21 399 27 405
rect 33 399 39 405
rect 45 399 51 405
rect 57 399 63 405
rect 69 399 75 405
rect 81 399 87 405
rect 93 399 99 405
rect 105 399 111 405
rect 117 399 123 405
rect 129 399 135 405
rect 141 399 147 405
rect 153 399 159 405
rect 165 399 171 405
rect 177 399 183 405
rect 189 399 195 405
rect 201 399 207 405
rect 213 399 219 405
rect 225 399 231 405
rect 237 399 243 405
rect 249 399 255 405
rect 261 399 267 405
rect 273 399 279 405
rect 285 399 291 405
rect 297 399 303 405
rect 309 399 315 405
rect 321 399 327 405
rect 333 399 339 405
rect 345 399 351 405
rect 357 399 363 405
rect 369 399 375 405
rect 381 399 387 405
rect 393 399 399 405
rect 405 399 411 405
rect 417 399 423 405
rect 429 399 435 405
rect 441 399 447 405
rect 453 399 459 405
rect 465 399 471 405
rect 477 399 483 405
rect 489 399 495 405
rect 501 399 507 405
rect 513 399 519 405
rect 525 399 531 405
rect 537 399 543 405
rect 549 399 555 405
rect 561 399 567 405
rect 573 399 579 405
rect 585 399 591 405
rect 597 399 603 405
rect 609 399 615 405
rect 621 399 627 405
rect 633 399 639 405
rect 645 399 651 405
rect 657 399 663 405
rect 669 399 675 405
rect 681 399 687 405
rect 693 399 699 405
rect 705 399 711 405
rect 717 399 723 405
rect 729 399 735 405
rect 741 399 747 405
rect 753 399 759 405
rect 765 399 771 405
rect 777 399 783 405
rect 789 399 795 405
rect 801 399 807 405
rect 813 399 819 405
rect 825 399 831 405
rect 837 399 843 405
rect 849 399 855 405
rect 861 399 867 405
rect 873 399 879 405
rect 885 399 891 405
rect 897 399 903 405
rect 909 399 915 405
rect 921 399 927 405
rect 933 399 939 405
rect 945 399 951 405
rect 957 399 963 405
rect 969 399 975 405
rect 981 399 987 405
rect 993 399 999 405
rect 1005 399 1011 405
rect 1017 399 1023 405
rect 1029 399 1035 405
rect 1041 399 1047 405
rect 1053 399 1059 405
rect 1065 399 1071 405
rect 1077 399 1083 405
rect 1089 399 1095 405
rect 1101 399 1107 405
rect 1113 399 1119 405
rect 1125 399 1131 405
rect 1137 399 1143 405
rect 1149 399 1155 405
rect 1161 399 1167 405
rect 1173 399 1179 405
rect 1185 399 1191 405
rect 1197 399 1203 405
rect 1209 399 1215 405
rect 1221 399 1227 405
rect 1233 399 1239 405
rect 1245 399 1251 405
rect 1257 399 1263 405
rect 1269 399 1275 405
rect 1281 399 1287 405
rect 1293 399 1299 405
rect 1305 399 1311 405
rect 1317 399 1323 405
rect 1329 399 1335 405
rect 1341 399 1347 405
rect 1353 399 1359 405
rect 1365 399 1371 405
rect 1377 399 1383 405
rect 1389 399 1395 405
rect 1401 399 1407 405
rect 1413 399 1419 405
rect 1425 399 1431 405
rect 1437 399 1443 405
rect 1449 399 1455 405
rect 1461 399 1467 405
rect 1473 399 1479 405
rect 1485 399 1491 405
rect 1497 399 1503 405
rect 1509 399 1512 405
rect -36 396 1512 399
rect -36 393 -24 396
rect -36 387 -33 393
rect -27 387 -24 393
rect -36 381 -24 387
rect -36 375 -33 381
rect -27 375 -24 381
rect -36 369 -24 375
rect -36 363 -33 369
rect -27 363 -24 369
rect -36 360 -24 363
rect 1500 393 1512 396
rect 1500 387 1503 393
rect 1509 387 1512 393
rect 1500 381 1512 387
rect 1500 375 1503 381
rect 1509 375 1512 381
rect 1500 369 1512 375
rect 1500 363 1503 369
rect 1509 363 1512 369
rect 1500 360 1512 363
rect -36 357 1512 360
rect -36 351 -33 357
rect -27 351 -21 357
rect -15 351 -9 357
rect -3 351 3 357
rect 9 351 15 357
rect 21 351 27 357
rect 33 351 39 357
rect 45 351 51 357
rect 57 351 63 357
rect 69 351 75 357
rect 81 351 87 357
rect 93 351 99 357
rect 105 351 111 357
rect 117 351 123 357
rect 129 351 135 357
rect 141 351 147 357
rect 153 351 159 357
rect 165 351 171 357
rect 177 351 183 357
rect 189 351 195 357
rect 201 351 207 357
rect 213 351 219 357
rect 225 351 231 357
rect 237 351 243 357
rect 249 351 255 357
rect 261 351 267 357
rect 273 351 279 357
rect 285 351 291 357
rect 297 351 303 357
rect 309 351 315 357
rect 321 351 327 357
rect 333 351 339 357
rect 345 351 351 357
rect 357 351 363 357
rect 369 351 375 357
rect 381 351 387 357
rect 393 351 399 357
rect 405 351 411 357
rect 417 351 423 357
rect 429 351 435 357
rect 441 351 447 357
rect 453 351 459 357
rect 465 351 471 357
rect 477 351 483 357
rect 489 351 495 357
rect 501 351 507 357
rect 513 351 519 357
rect 525 351 531 357
rect 537 351 543 357
rect 549 351 555 357
rect 561 351 567 357
rect 573 351 579 357
rect 585 351 591 357
rect 597 351 603 357
rect 609 351 615 357
rect 621 351 627 357
rect 633 351 639 357
rect 645 351 651 357
rect 657 351 663 357
rect 669 351 675 357
rect 681 351 687 357
rect 693 351 699 357
rect 705 351 711 357
rect 717 351 723 357
rect 729 351 735 357
rect 741 351 747 357
rect 753 351 759 357
rect 765 351 771 357
rect 777 351 783 357
rect 789 351 795 357
rect 801 351 807 357
rect 813 351 819 357
rect 825 351 831 357
rect 837 351 843 357
rect 849 351 855 357
rect 861 351 867 357
rect 873 351 879 357
rect 885 351 891 357
rect 897 351 903 357
rect 909 351 915 357
rect 921 351 927 357
rect 933 351 939 357
rect 945 351 951 357
rect 957 351 963 357
rect 969 351 975 357
rect 981 351 987 357
rect 993 351 999 357
rect 1005 351 1011 357
rect 1017 351 1023 357
rect 1029 351 1035 357
rect 1041 351 1047 357
rect 1053 351 1059 357
rect 1065 351 1071 357
rect 1077 351 1083 357
rect 1089 351 1095 357
rect 1101 351 1107 357
rect 1113 351 1119 357
rect 1125 351 1131 357
rect 1137 351 1143 357
rect 1149 351 1155 357
rect 1161 351 1167 357
rect 1173 351 1179 357
rect 1185 351 1191 357
rect 1197 351 1203 357
rect 1209 351 1215 357
rect 1221 351 1227 357
rect 1233 351 1239 357
rect 1245 351 1251 357
rect 1257 351 1263 357
rect 1269 351 1275 357
rect 1281 351 1287 357
rect 1293 351 1299 357
rect 1305 351 1311 357
rect 1317 351 1323 357
rect 1329 351 1335 357
rect 1341 351 1347 357
rect 1353 351 1359 357
rect 1365 351 1371 357
rect 1377 351 1383 357
rect 1389 351 1395 357
rect 1401 351 1407 357
rect 1413 351 1419 357
rect 1425 351 1431 357
rect 1437 351 1443 357
rect 1449 351 1455 357
rect 1461 351 1467 357
rect 1473 351 1479 357
rect 1485 351 1491 357
rect 1497 351 1503 357
rect 1509 351 1512 357
rect -36 348 1512 351
rect 1524 597 1536 603
rect 1524 591 1527 597
rect 1533 591 1536 597
rect 1524 585 1536 591
rect 1524 579 1527 585
rect 1533 579 1536 585
rect 1524 573 1536 579
rect 1524 567 1527 573
rect 1533 567 1536 573
rect 1524 561 1536 567
rect 1524 555 1527 561
rect 1533 555 1536 561
rect 1524 549 1536 555
rect 1524 543 1527 549
rect 1533 543 1536 549
rect 1524 537 1536 543
rect 1524 531 1527 537
rect 1533 531 1536 537
rect 1524 525 1536 531
rect 1524 519 1527 525
rect 1533 519 1536 525
rect 1524 513 1536 519
rect 1524 507 1527 513
rect 1533 507 1536 513
rect 1524 501 1536 507
rect 1524 495 1527 501
rect 1533 495 1536 501
rect 1524 489 1536 495
rect 1524 483 1527 489
rect 1533 483 1536 489
rect 1524 477 1536 483
rect 1524 471 1527 477
rect 1533 471 1536 477
rect 1524 465 1536 471
rect 1524 459 1527 465
rect 1533 459 1536 465
rect 1524 453 1536 459
rect 1524 447 1527 453
rect 1533 447 1536 453
rect 1524 441 1536 447
rect 1524 435 1527 441
rect 1533 435 1536 441
rect 1524 429 1536 435
rect 1524 423 1527 429
rect 1533 423 1536 429
rect 1524 417 1536 423
rect 1524 411 1527 417
rect 1533 411 1536 417
rect 1524 405 1536 411
rect 1524 399 1527 405
rect 1533 399 1536 405
rect 1524 393 1536 399
rect 1524 387 1527 393
rect 1533 387 1536 393
rect 1524 381 1536 387
rect 1524 375 1527 381
rect 1533 375 1536 381
rect 1524 369 1536 375
rect 1524 363 1527 369
rect 1533 363 1536 369
rect 1524 357 1536 363
rect 1524 351 1527 357
rect 1533 351 1536 357
rect -60 339 -57 345
rect -51 339 -48 345
rect -60 336 -48 339
rect 1524 345 1536 351
rect 1524 339 1527 345
rect 1533 339 1536 345
rect 1524 336 1536 339
rect -60 333 1536 336
rect -60 327 -57 333
rect -51 327 -45 333
rect -39 327 -33 333
rect -27 327 -21 333
rect -15 327 -9 333
rect -3 327 3 333
rect 9 327 15 333
rect 21 327 27 333
rect 33 327 39 333
rect 45 327 51 333
rect 57 327 63 333
rect 69 327 75 333
rect 81 327 87 333
rect 93 327 99 333
rect 105 327 111 333
rect 117 327 123 333
rect 129 327 135 333
rect 141 327 147 333
rect 153 327 159 333
rect 165 327 171 333
rect 177 327 183 333
rect 189 327 195 333
rect 201 327 207 333
rect 213 327 219 333
rect 225 327 231 333
rect 237 327 243 333
rect 249 327 255 333
rect 261 327 267 333
rect 273 327 279 333
rect 285 327 291 333
rect 297 327 303 333
rect 309 327 315 333
rect 321 327 327 333
rect 333 327 339 333
rect 345 327 351 333
rect 357 327 363 333
rect 369 327 375 333
rect 381 327 387 333
rect 393 327 399 333
rect 405 327 411 333
rect 417 327 423 333
rect 429 327 435 333
rect 441 327 447 333
rect 453 327 459 333
rect 465 327 471 333
rect 477 327 483 333
rect 489 327 495 333
rect 501 327 507 333
rect 513 327 519 333
rect 525 327 531 333
rect 537 327 543 333
rect 549 327 555 333
rect 561 327 567 333
rect 573 327 579 333
rect 585 327 591 333
rect 597 327 603 333
rect 609 327 615 333
rect 621 327 627 333
rect 633 327 639 333
rect 645 327 651 333
rect 657 327 663 333
rect 669 327 675 333
rect 681 327 687 333
rect 693 327 699 333
rect 705 327 711 333
rect 717 327 723 333
rect 729 327 735 333
rect 741 327 747 333
rect 753 327 759 333
rect 765 327 771 333
rect 777 327 783 333
rect 789 327 795 333
rect 801 327 807 333
rect 813 327 819 333
rect 825 327 831 333
rect 837 327 843 333
rect 849 327 855 333
rect 861 327 867 333
rect 873 327 879 333
rect 885 327 891 333
rect 897 327 903 333
rect 909 327 915 333
rect 921 327 927 333
rect 933 327 939 333
rect 945 327 951 333
rect 957 327 963 333
rect 969 327 975 333
rect 981 327 987 333
rect 993 327 999 333
rect 1005 327 1011 333
rect 1017 327 1023 333
rect 1029 327 1035 333
rect 1041 327 1047 333
rect 1053 327 1059 333
rect 1065 327 1071 333
rect 1077 327 1083 333
rect 1089 327 1095 333
rect 1101 327 1107 333
rect 1113 327 1119 333
rect 1125 327 1131 333
rect 1137 327 1143 333
rect 1149 327 1155 333
rect 1161 327 1167 333
rect 1173 327 1179 333
rect 1185 327 1191 333
rect 1197 327 1203 333
rect 1209 327 1215 333
rect 1221 327 1227 333
rect 1233 327 1239 333
rect 1245 327 1251 333
rect 1257 327 1263 333
rect 1269 327 1275 333
rect 1281 327 1287 333
rect 1293 327 1299 333
rect 1305 327 1311 333
rect 1317 327 1323 333
rect 1329 327 1335 333
rect 1341 327 1347 333
rect 1353 327 1359 333
rect 1365 327 1371 333
rect 1377 327 1383 333
rect 1389 327 1395 333
rect 1401 327 1407 333
rect 1413 327 1419 333
rect 1425 327 1431 333
rect 1437 327 1443 333
rect 1449 327 1455 333
rect 1461 327 1467 333
rect 1473 327 1479 333
rect 1485 327 1491 333
rect 1497 327 1503 333
rect 1509 327 1515 333
rect 1521 327 1527 333
rect 1533 327 1536 333
rect -60 324 1536 327
rect -60 321 -48 324
rect -60 315 -57 321
rect -51 315 -48 321
rect -60 309 -48 315
rect 1524 321 1536 324
rect 1524 315 1527 321
rect 1533 315 1536 321
rect -60 303 -57 309
rect -51 303 -48 309
rect -60 297 -48 303
rect -12 309 192 312
rect -12 303 -9 309
rect -3 303 3 309
rect 9 303 15 309
rect 21 303 27 309
rect 33 303 39 309
rect 45 303 51 309
rect 57 303 63 309
rect 69 303 75 309
rect 81 303 87 309
rect 93 303 99 309
rect 105 303 111 309
rect 117 303 123 309
rect 129 303 135 309
rect 141 303 147 309
rect 153 303 159 309
rect 165 303 171 309
rect 177 303 183 309
rect 189 303 192 309
rect -12 300 192 303
rect 216 309 252 312
rect 216 303 219 309
rect 225 303 231 309
rect 237 303 243 309
rect 249 303 252 309
rect 216 300 252 303
rect 264 309 300 312
rect 264 303 267 309
rect 273 303 279 309
rect 285 303 291 309
rect 297 303 300 309
rect 264 300 300 303
rect 312 309 348 312
rect 312 303 315 309
rect 321 303 327 309
rect 333 303 339 309
rect 345 303 348 309
rect 312 300 348 303
rect 360 309 396 312
rect 360 303 363 309
rect 369 303 375 309
rect 381 303 387 309
rect 393 303 396 309
rect 360 300 396 303
rect 432 309 468 312
rect 432 303 435 309
rect 441 303 447 309
rect 453 303 459 309
rect 465 303 468 309
rect 432 300 468 303
rect 480 309 516 312
rect 480 303 483 309
rect 489 303 495 309
rect 501 303 507 309
rect 513 303 516 309
rect 480 300 516 303
rect 528 309 564 312
rect 528 303 531 309
rect 537 303 543 309
rect 549 303 555 309
rect 561 303 564 309
rect 528 300 564 303
rect 576 309 612 312
rect 576 303 579 309
rect 585 303 591 309
rect 597 303 603 309
rect 609 303 612 309
rect 576 300 612 303
rect 648 309 684 312
rect 648 303 651 309
rect 657 303 663 309
rect 669 303 675 309
rect 681 303 684 309
rect 648 300 684 303
rect 696 309 732 312
rect 696 303 699 309
rect 705 303 711 309
rect 717 303 723 309
rect 729 303 732 309
rect 696 300 732 303
rect 744 309 780 312
rect 744 303 747 309
rect 753 303 759 309
rect 765 303 771 309
rect 777 303 780 309
rect 744 300 780 303
rect 792 309 828 312
rect 792 303 795 309
rect 801 303 807 309
rect 813 303 819 309
rect 825 303 828 309
rect 792 300 828 303
rect 864 309 876 312
rect 864 303 867 309
rect 873 303 876 309
rect 864 300 876 303
rect 912 309 948 312
rect 912 303 915 309
rect 921 303 927 309
rect 933 303 939 309
rect 945 303 948 309
rect 912 300 948 303
rect 960 309 996 312
rect 960 303 963 309
rect 969 303 975 309
rect 981 303 987 309
rect 993 303 996 309
rect 960 300 996 303
rect 1008 309 1044 312
rect 1008 303 1011 309
rect 1017 303 1023 309
rect 1029 303 1035 309
rect 1041 303 1044 309
rect 1008 300 1044 303
rect 1080 309 1116 312
rect 1080 303 1083 309
rect 1089 303 1095 309
rect 1101 303 1107 309
rect 1113 303 1116 309
rect 1080 300 1116 303
rect 1128 309 1164 312
rect 1128 303 1131 309
rect 1137 303 1143 309
rect 1149 303 1155 309
rect 1161 303 1164 309
rect 1128 300 1164 303
rect 1176 309 1212 312
rect 1176 303 1179 309
rect 1185 303 1191 309
rect 1197 303 1203 309
rect 1209 303 1212 309
rect 1176 300 1212 303
rect 1224 309 1260 312
rect 1224 303 1227 309
rect 1233 303 1239 309
rect 1245 303 1251 309
rect 1257 303 1260 309
rect 1224 300 1260 303
rect 1296 309 1332 312
rect 1296 303 1299 309
rect 1305 303 1311 309
rect 1317 303 1323 309
rect 1329 303 1332 309
rect 1296 300 1332 303
rect 1344 309 1380 312
rect 1344 303 1347 309
rect 1353 303 1359 309
rect 1365 303 1371 309
rect 1377 303 1380 309
rect 1344 300 1380 303
rect 1392 309 1428 312
rect 1392 303 1395 309
rect 1401 303 1407 309
rect 1413 303 1419 309
rect 1425 303 1428 309
rect 1392 300 1428 303
rect 1440 309 1476 312
rect 1440 303 1443 309
rect 1449 303 1455 309
rect 1461 303 1467 309
rect 1473 303 1476 309
rect 1440 300 1476 303
rect 1524 309 1536 315
rect 1524 303 1527 309
rect 1533 303 1536 309
rect -60 291 -57 297
rect -51 291 -48 297
rect -60 285 -48 291
rect -60 279 -57 285
rect -51 279 -48 285
rect -60 273 -48 279
rect -60 267 -57 273
rect -51 267 -48 273
rect -60 261 -48 267
rect -60 255 -57 261
rect -51 255 -48 261
rect -60 249 -48 255
rect -12 285 0 288
rect -12 279 -9 285
rect -3 279 0 285
rect -12 273 0 279
rect -12 267 -9 273
rect -3 267 0 273
rect -12 261 0 267
rect -12 255 -9 261
rect -3 255 0 261
rect -12 252 0 255
rect 12 285 24 300
rect 12 279 15 285
rect 21 279 24 285
rect 12 273 24 279
rect 12 267 15 273
rect 21 267 24 273
rect 12 261 24 267
rect 12 255 15 261
rect 21 255 24 261
rect 12 252 24 255
rect 36 285 48 288
rect 36 279 39 285
rect 45 279 48 285
rect 36 273 48 279
rect 36 267 39 273
rect 45 267 48 273
rect 36 261 48 267
rect 36 255 39 261
rect 45 255 48 261
rect 36 252 48 255
rect 60 285 72 300
rect 60 279 63 285
rect 69 279 72 285
rect 60 273 72 279
rect 60 267 63 273
rect 69 267 72 273
rect 60 261 72 267
rect 60 255 63 261
rect 69 255 72 261
rect 60 252 72 255
rect 84 285 96 288
rect 84 279 87 285
rect 93 279 96 285
rect 84 273 96 279
rect 84 267 87 273
rect 93 267 96 273
rect 84 261 96 267
rect 84 255 87 261
rect 93 255 96 261
rect 84 252 96 255
rect 108 285 120 300
rect 108 279 111 285
rect 117 279 120 285
rect 108 273 120 279
rect 108 267 111 273
rect 117 267 120 273
rect 108 261 120 267
rect 108 255 111 261
rect 117 255 120 261
rect 108 252 120 255
rect 132 285 144 288
rect 132 279 135 285
rect 141 279 144 285
rect 132 273 144 279
rect 132 267 135 273
rect 141 267 144 273
rect 132 261 144 267
rect 132 255 135 261
rect 141 255 144 261
rect 132 252 144 255
rect 156 285 168 300
rect 1524 297 1536 303
rect 1524 291 1527 297
rect 1533 291 1536 297
rect 156 279 159 285
rect 165 279 168 285
rect 156 273 168 279
rect 156 267 159 273
rect 165 267 168 273
rect 156 261 168 267
rect 156 255 159 261
rect 165 255 168 261
rect 156 252 168 255
rect 180 285 192 288
rect 180 279 183 285
rect 189 279 192 285
rect 180 273 192 279
rect 180 267 183 273
rect 189 267 192 273
rect 180 261 192 267
rect 180 255 183 261
rect 189 255 192 261
rect 180 252 192 255
rect 204 285 216 288
rect 204 279 207 285
rect 213 279 216 285
rect 204 273 216 279
rect 204 267 207 273
rect 213 267 216 273
rect 204 261 216 267
rect 204 255 207 261
rect 213 255 216 261
rect 204 252 216 255
rect 300 285 312 288
rect 300 279 303 285
rect 309 279 312 285
rect 300 273 312 279
rect 300 267 303 273
rect 309 267 312 273
rect 300 261 312 267
rect 300 255 303 261
rect 309 255 312 261
rect 300 252 312 255
rect 396 285 408 288
rect 396 279 399 285
rect 405 279 408 285
rect 396 273 408 279
rect 396 267 399 273
rect 405 267 408 273
rect 396 261 408 267
rect 396 255 399 261
rect 405 255 408 261
rect 396 252 408 255
rect 420 285 432 288
rect 420 279 423 285
rect 429 279 432 285
rect 420 273 432 279
rect 420 267 423 273
rect 429 267 432 273
rect 420 261 432 267
rect 420 255 423 261
rect 429 255 432 261
rect 420 252 432 255
rect 516 285 528 288
rect 516 279 519 285
rect 525 279 528 285
rect 516 273 528 279
rect 516 267 519 273
rect 525 267 528 273
rect 516 261 528 267
rect 516 255 519 261
rect 525 255 528 261
rect 516 252 528 255
rect 612 285 624 288
rect 612 279 615 285
rect 621 279 624 285
rect 612 273 624 279
rect 612 267 615 273
rect 621 267 624 273
rect 612 261 624 267
rect 612 255 615 261
rect 621 255 624 261
rect 612 252 624 255
rect 636 285 648 288
rect 636 279 639 285
rect 645 279 648 285
rect 636 273 648 279
rect 636 267 639 273
rect 645 267 648 273
rect 636 261 648 267
rect 636 255 639 261
rect 645 255 648 261
rect 636 252 648 255
rect 732 285 744 288
rect 732 279 735 285
rect 741 279 744 285
rect 732 273 744 279
rect 732 267 735 273
rect 741 267 744 273
rect 732 261 744 267
rect 732 255 735 261
rect 741 255 744 261
rect 732 252 744 255
rect 828 285 840 288
rect 828 279 831 285
rect 837 279 840 285
rect 828 273 840 279
rect 828 267 831 273
rect 837 267 840 273
rect 828 261 840 267
rect 828 255 831 261
rect 837 255 840 261
rect 828 252 840 255
rect 852 285 864 288
rect 852 279 855 285
rect 861 279 864 285
rect 852 273 864 279
rect 852 267 855 273
rect 861 267 864 273
rect 852 261 864 267
rect 852 255 855 261
rect 861 255 864 261
rect 852 252 864 255
rect 876 285 888 288
rect 876 279 879 285
rect 885 279 888 285
rect 876 273 888 279
rect 876 267 879 273
rect 885 267 888 273
rect 876 261 888 267
rect 876 255 879 261
rect 885 255 888 261
rect 876 252 888 255
rect 900 285 912 288
rect 900 279 903 285
rect 909 279 912 285
rect 900 273 912 279
rect 900 267 903 273
rect 909 267 912 273
rect 900 261 912 267
rect 900 255 903 261
rect 909 255 912 261
rect 900 252 912 255
rect 1044 285 1056 288
rect 1044 279 1047 285
rect 1053 279 1056 285
rect 1044 273 1056 279
rect 1044 267 1047 273
rect 1053 267 1056 273
rect 1044 261 1056 267
rect 1044 255 1047 261
rect 1053 255 1056 261
rect 1044 252 1056 255
rect 1068 285 1080 288
rect 1068 279 1071 285
rect 1077 279 1080 285
rect 1068 273 1080 279
rect 1068 267 1071 273
rect 1077 267 1080 273
rect 1068 261 1080 267
rect 1068 255 1071 261
rect 1077 255 1080 261
rect 1068 252 1080 255
rect 1092 285 1104 288
rect 1092 279 1095 285
rect 1101 279 1104 285
rect 1092 273 1104 279
rect 1092 267 1095 273
rect 1101 267 1104 273
rect 1092 261 1104 267
rect 1092 255 1095 261
rect 1101 255 1104 261
rect 1092 252 1104 255
rect 1116 285 1128 288
rect 1116 279 1119 285
rect 1125 279 1128 285
rect 1116 273 1128 279
rect 1116 267 1119 273
rect 1125 267 1128 273
rect 1116 261 1128 267
rect 1116 255 1119 261
rect 1125 255 1128 261
rect 1116 252 1128 255
rect 1140 285 1152 288
rect 1140 279 1143 285
rect 1149 279 1152 285
rect 1140 273 1152 279
rect 1140 267 1143 273
rect 1149 267 1152 273
rect 1140 261 1152 267
rect 1140 255 1143 261
rect 1149 255 1152 261
rect 1140 252 1152 255
rect 1164 285 1176 288
rect 1164 279 1167 285
rect 1173 279 1176 285
rect 1164 273 1176 279
rect 1164 267 1167 273
rect 1173 267 1176 273
rect 1164 261 1176 267
rect 1164 255 1167 261
rect 1173 255 1176 261
rect 1164 252 1176 255
rect 1188 285 1200 288
rect 1188 279 1191 285
rect 1197 279 1200 285
rect 1188 273 1200 279
rect 1188 267 1191 273
rect 1197 267 1200 273
rect 1188 261 1200 267
rect 1188 255 1191 261
rect 1197 255 1200 261
rect 1188 252 1200 255
rect 1212 285 1224 288
rect 1212 279 1215 285
rect 1221 279 1224 285
rect 1212 273 1224 279
rect 1212 267 1215 273
rect 1221 267 1224 273
rect 1212 261 1224 267
rect 1212 255 1215 261
rect 1221 255 1224 261
rect 1212 252 1224 255
rect 1236 285 1248 288
rect 1236 279 1239 285
rect 1245 279 1248 285
rect 1236 273 1248 279
rect 1236 267 1239 273
rect 1245 267 1248 273
rect 1236 261 1248 267
rect 1236 255 1239 261
rect 1245 255 1248 261
rect 1236 252 1248 255
rect 1260 285 1272 288
rect 1260 279 1263 285
rect 1269 279 1272 285
rect 1260 273 1272 279
rect 1260 267 1263 273
rect 1269 267 1272 273
rect 1260 261 1272 267
rect 1260 255 1263 261
rect 1269 255 1272 261
rect 1260 252 1272 255
rect 1284 285 1296 288
rect 1284 279 1287 285
rect 1293 279 1296 285
rect 1284 273 1296 279
rect 1284 267 1287 273
rect 1293 267 1296 273
rect 1284 261 1296 267
rect 1284 255 1287 261
rect 1293 255 1296 261
rect 1284 252 1296 255
rect 1308 285 1320 288
rect 1308 279 1311 285
rect 1317 279 1320 285
rect 1308 273 1320 279
rect 1308 267 1311 273
rect 1317 267 1320 273
rect 1308 261 1320 267
rect 1308 255 1311 261
rect 1317 255 1320 261
rect 1308 252 1320 255
rect 1332 285 1344 288
rect 1332 279 1335 285
rect 1341 279 1344 285
rect 1332 273 1344 279
rect 1332 267 1335 273
rect 1341 267 1344 273
rect 1332 261 1344 267
rect 1332 255 1335 261
rect 1341 255 1344 261
rect 1332 252 1344 255
rect 1356 285 1368 288
rect 1356 279 1359 285
rect 1365 279 1368 285
rect 1356 273 1368 279
rect 1356 267 1359 273
rect 1365 267 1368 273
rect 1356 261 1368 267
rect 1356 255 1359 261
rect 1365 255 1368 261
rect 1356 252 1368 255
rect 1380 285 1392 288
rect 1380 279 1383 285
rect 1389 279 1392 285
rect 1380 273 1392 279
rect 1380 267 1383 273
rect 1389 267 1392 273
rect 1380 261 1392 267
rect 1380 255 1383 261
rect 1389 255 1392 261
rect 1380 252 1392 255
rect 1404 285 1416 288
rect 1404 279 1407 285
rect 1413 279 1416 285
rect 1404 273 1416 279
rect 1404 267 1407 273
rect 1413 267 1416 273
rect 1404 261 1416 267
rect 1404 255 1407 261
rect 1413 255 1416 261
rect 1404 252 1416 255
rect 1428 285 1440 288
rect 1428 279 1431 285
rect 1437 279 1440 285
rect 1428 273 1440 279
rect 1428 267 1431 273
rect 1437 267 1440 273
rect 1428 261 1440 267
rect 1428 255 1431 261
rect 1437 255 1440 261
rect 1428 252 1440 255
rect 1452 285 1464 288
rect 1452 279 1455 285
rect 1461 279 1464 285
rect 1452 273 1464 279
rect 1452 267 1455 273
rect 1461 267 1464 273
rect 1452 261 1464 267
rect 1452 255 1455 261
rect 1461 255 1464 261
rect 1452 252 1464 255
rect 1476 285 1488 288
rect 1476 279 1479 285
rect 1485 279 1488 285
rect 1476 273 1488 279
rect 1476 267 1479 273
rect 1485 267 1488 273
rect 1476 261 1488 267
rect 1476 255 1479 261
rect 1485 255 1488 261
rect 1476 252 1488 255
rect 1524 285 1536 291
rect 1524 279 1527 285
rect 1533 279 1536 285
rect 1524 273 1536 279
rect 1524 267 1527 273
rect 1533 267 1536 273
rect 1524 261 1536 267
rect 1524 255 1527 261
rect 1533 255 1536 261
rect -60 243 -57 249
rect -51 243 -48 249
rect -60 237 -48 243
rect -60 231 -57 237
rect -51 231 -48 237
rect -60 225 -48 231
rect -60 219 -57 225
rect -51 219 -48 225
rect -60 216 -48 219
rect 1524 249 1536 255
rect 1524 243 1527 249
rect 1533 243 1536 249
rect 1524 237 1536 243
rect 1524 231 1527 237
rect 1533 231 1536 237
rect 1524 225 1536 231
rect 1524 219 1527 225
rect 1533 219 1536 225
rect 1524 216 1536 219
rect -60 213 1536 216
rect -60 207 -57 213
rect -51 207 -45 213
rect -39 207 -33 213
rect -27 207 -21 213
rect -15 207 -9 213
rect -3 207 3 213
rect 9 207 15 213
rect 21 207 27 213
rect 33 207 39 213
rect 45 207 51 213
rect 57 207 63 213
rect 69 207 75 213
rect 81 207 87 213
rect 93 207 99 213
rect 105 207 111 213
rect 117 207 123 213
rect 129 207 135 213
rect 141 207 147 213
rect 153 207 159 213
rect 165 207 171 213
rect 177 207 183 213
rect 189 207 195 213
rect 201 207 207 213
rect 213 207 219 213
rect 225 207 231 213
rect 237 207 243 213
rect 249 207 255 213
rect 261 207 267 213
rect 273 207 279 213
rect 285 207 291 213
rect 297 207 303 213
rect 309 207 315 213
rect 321 207 327 213
rect 333 207 339 213
rect 345 207 351 213
rect 357 207 363 213
rect 369 207 375 213
rect 381 207 387 213
rect 393 207 399 213
rect 405 207 411 213
rect 417 207 423 213
rect 429 207 435 213
rect 441 207 447 213
rect 453 207 459 213
rect 465 207 471 213
rect 477 207 483 213
rect 489 207 495 213
rect 501 207 507 213
rect 513 207 519 213
rect 525 207 531 213
rect 537 207 543 213
rect 549 207 555 213
rect 561 207 567 213
rect 573 207 579 213
rect 585 207 591 213
rect 597 207 603 213
rect 609 207 615 213
rect 621 207 627 213
rect 633 207 639 213
rect 645 207 651 213
rect 657 207 663 213
rect 669 207 675 213
rect 681 207 687 213
rect 693 207 699 213
rect 705 207 711 213
rect 717 207 723 213
rect 729 207 735 213
rect 741 207 747 213
rect 753 207 759 213
rect 765 207 771 213
rect 777 207 783 213
rect 789 207 795 213
rect 801 207 807 213
rect 813 207 819 213
rect 825 207 831 213
rect 837 207 843 213
rect 849 207 855 213
rect 861 207 867 213
rect 873 207 879 213
rect 885 207 891 213
rect 897 207 903 213
rect 909 207 915 213
rect 921 207 927 213
rect 933 207 939 213
rect 945 207 951 213
rect 957 207 963 213
rect 969 207 975 213
rect 981 207 987 213
rect 993 207 999 213
rect 1005 207 1011 213
rect 1017 207 1023 213
rect 1029 207 1035 213
rect 1041 207 1047 213
rect 1053 207 1059 213
rect 1065 207 1071 213
rect 1077 207 1083 213
rect 1089 207 1095 213
rect 1101 207 1107 213
rect 1113 207 1119 213
rect 1125 207 1131 213
rect 1137 207 1143 213
rect 1149 207 1155 213
rect 1161 207 1167 213
rect 1173 207 1179 213
rect 1185 207 1191 213
rect 1197 207 1203 213
rect 1209 207 1215 213
rect 1221 207 1227 213
rect 1233 207 1239 213
rect 1245 207 1251 213
rect 1257 207 1263 213
rect 1269 207 1275 213
rect 1281 207 1287 213
rect 1293 207 1299 213
rect 1305 207 1311 213
rect 1317 207 1323 213
rect 1329 207 1335 213
rect 1341 207 1347 213
rect 1353 207 1359 213
rect 1365 207 1371 213
rect 1377 207 1383 213
rect 1389 207 1395 213
rect 1401 207 1407 213
rect 1413 207 1419 213
rect 1425 207 1431 213
rect 1437 207 1443 213
rect 1449 207 1455 213
rect 1461 207 1467 213
rect 1473 207 1479 213
rect 1485 207 1491 213
rect 1497 207 1503 213
rect 1509 207 1515 213
rect 1521 207 1527 213
rect 1533 207 1536 213
rect -60 204 1536 207
rect -60 201 -48 204
rect -60 195 -57 201
rect -51 195 -48 201
rect -60 189 -48 195
rect -60 183 -57 189
rect -51 183 -48 189
rect -60 177 -48 183
rect -60 171 -57 177
rect -51 171 -48 177
rect -60 165 -48 171
rect -60 159 -57 165
rect -51 159 -48 165
rect -60 153 -48 159
rect -60 147 -57 153
rect -51 147 -48 153
rect -60 141 -48 147
rect -60 135 -57 141
rect -51 135 -48 141
rect -60 129 -48 135
rect -60 123 -57 129
rect -51 123 -48 129
rect -60 117 -48 123
rect -60 111 -57 117
rect -51 111 -48 117
rect -60 105 -48 111
rect -60 99 -57 105
rect -51 99 -48 105
rect -60 96 -48 99
rect 1524 201 1536 204
rect 1524 195 1527 201
rect 1533 195 1536 201
rect 1524 189 1536 195
rect 1524 183 1527 189
rect 1533 183 1536 189
rect 1524 177 1536 183
rect 1524 171 1527 177
rect 1533 171 1536 177
rect 1524 165 1536 171
rect 1524 159 1527 165
rect 1533 159 1536 165
rect 1524 153 1536 159
rect 1524 147 1527 153
rect 1533 147 1536 153
rect 1524 141 1536 147
rect 1524 135 1527 141
rect 1533 135 1536 141
rect 1524 129 1536 135
rect 1524 123 1527 129
rect 1533 123 1536 129
rect 1524 117 1536 123
rect 1524 111 1527 117
rect 1533 111 1536 117
rect 1524 105 1536 111
rect 1524 99 1527 105
rect 1533 99 1536 105
rect 1524 96 1536 99
rect -60 93 1536 96
rect -60 87 -57 93
rect -51 87 -45 93
rect -39 87 -33 93
rect -27 87 -21 93
rect -15 87 -9 93
rect -3 87 3 93
rect 9 87 15 93
rect 21 87 27 93
rect 33 87 39 93
rect 45 87 51 93
rect 57 87 63 93
rect 69 87 75 93
rect 81 87 87 93
rect 93 87 99 93
rect 105 87 111 93
rect 117 87 123 93
rect 129 87 135 93
rect 141 87 147 93
rect 153 87 159 93
rect 165 87 171 93
rect 177 87 183 93
rect 189 87 195 93
rect 201 87 207 93
rect 213 87 219 93
rect 225 87 231 93
rect 237 87 243 93
rect 249 87 255 93
rect 261 87 267 93
rect 273 87 279 93
rect 285 87 291 93
rect 297 87 303 93
rect 309 87 315 93
rect 321 87 327 93
rect 333 87 339 93
rect 345 87 351 93
rect 357 87 363 93
rect 369 87 375 93
rect 381 87 387 93
rect 393 87 399 93
rect 405 87 411 93
rect 417 87 423 93
rect 429 87 435 93
rect 441 87 447 93
rect 453 87 459 93
rect 465 87 471 93
rect 477 87 483 93
rect 489 87 495 93
rect 501 87 507 93
rect 513 87 519 93
rect 525 87 531 93
rect 537 87 543 93
rect 549 87 555 93
rect 561 87 567 93
rect 573 87 579 93
rect 585 87 591 93
rect 597 87 603 93
rect 609 87 615 93
rect 621 87 627 93
rect 633 87 639 93
rect 645 87 651 93
rect 657 87 663 93
rect 669 87 675 93
rect 681 87 687 93
rect 693 87 699 93
rect 705 87 711 93
rect 717 87 723 93
rect 729 87 735 93
rect 741 87 747 93
rect 753 87 759 93
rect 765 87 771 93
rect 777 87 783 93
rect 789 87 795 93
rect 801 87 807 93
rect 813 87 819 93
rect 825 87 831 93
rect 837 87 843 93
rect 849 87 855 93
rect 861 87 867 93
rect 873 87 879 93
rect 885 87 891 93
rect 897 87 903 93
rect 909 87 915 93
rect 921 87 927 93
rect 933 87 939 93
rect 945 87 951 93
rect 957 87 963 93
rect 969 87 975 93
rect 981 87 987 93
rect 993 87 999 93
rect 1005 87 1011 93
rect 1017 87 1023 93
rect 1029 87 1035 93
rect 1041 87 1047 93
rect 1053 87 1059 93
rect 1065 87 1071 93
rect 1077 87 1083 93
rect 1089 87 1095 93
rect 1101 87 1107 93
rect 1113 87 1119 93
rect 1125 87 1131 93
rect 1137 87 1143 93
rect 1149 87 1155 93
rect 1161 87 1167 93
rect 1173 87 1179 93
rect 1185 87 1191 93
rect 1197 87 1203 93
rect 1209 87 1215 93
rect 1221 87 1227 93
rect 1233 87 1239 93
rect 1245 87 1251 93
rect 1257 87 1263 93
rect 1269 87 1275 93
rect 1281 87 1287 93
rect 1293 87 1299 93
rect 1305 87 1311 93
rect 1317 87 1323 93
rect 1329 87 1335 93
rect 1341 87 1347 93
rect 1353 87 1359 93
rect 1365 87 1371 93
rect 1377 87 1383 93
rect 1389 87 1395 93
rect 1401 87 1407 93
rect 1413 87 1419 93
rect 1425 87 1431 93
rect 1437 87 1443 93
rect 1449 87 1455 93
rect 1461 87 1467 93
rect 1473 87 1479 93
rect 1485 87 1491 93
rect 1497 87 1503 93
rect 1509 87 1515 93
rect 1521 87 1527 93
rect 1533 87 1536 93
rect -60 84 1536 87
rect -60 81 -48 84
rect -60 75 -57 81
rect -51 75 -48 81
rect -60 69 -48 75
rect 1524 81 1536 84
rect 1524 75 1527 81
rect 1533 75 1536 81
rect -60 63 -57 69
rect -51 63 -48 69
rect -60 57 -48 63
rect 0 69 36 72
rect 0 63 3 69
rect 9 63 15 69
rect 21 63 27 69
rect 33 63 36 69
rect 0 60 36 63
rect 48 69 84 72
rect 48 63 51 69
rect 57 63 63 69
rect 69 63 75 69
rect 81 63 84 69
rect 48 60 84 63
rect 96 69 132 72
rect 96 63 99 69
rect 105 63 111 69
rect 117 63 123 69
rect 129 63 132 69
rect 96 60 132 63
rect 144 69 180 72
rect 144 63 147 69
rect 153 63 159 69
rect 165 63 171 69
rect 177 63 180 69
rect 144 60 180 63
rect 216 69 252 72
rect 216 63 219 69
rect 225 63 231 69
rect 237 63 243 69
rect 249 63 252 69
rect 216 60 252 63
rect 264 69 300 72
rect 264 63 267 69
rect 273 63 279 69
rect 285 63 291 69
rect 297 63 300 69
rect 264 60 300 63
rect 312 69 348 72
rect 312 63 315 69
rect 321 63 327 69
rect 333 63 339 69
rect 345 63 348 69
rect 312 60 348 63
rect 360 69 396 72
rect 360 63 363 69
rect 369 63 375 69
rect 381 63 387 69
rect 393 63 396 69
rect 360 60 396 63
rect 432 69 468 72
rect 432 63 435 69
rect 441 63 447 69
rect 453 63 459 69
rect 465 63 468 69
rect 432 60 468 63
rect 480 69 516 72
rect 480 63 483 69
rect 489 63 495 69
rect 501 63 507 69
rect 513 63 516 69
rect 480 60 516 63
rect 528 69 564 72
rect 528 63 531 69
rect 537 63 543 69
rect 549 63 555 69
rect 561 63 564 69
rect 528 60 564 63
rect 576 69 612 72
rect 576 63 579 69
rect 585 63 591 69
rect 597 63 603 69
rect 609 63 612 69
rect 576 60 612 63
rect 648 69 684 72
rect 648 63 651 69
rect 657 63 663 69
rect 669 63 675 69
rect 681 63 684 69
rect 648 60 684 63
rect 696 69 732 72
rect 696 63 699 69
rect 705 63 711 69
rect 717 63 723 69
rect 729 63 732 69
rect 696 60 732 63
rect 744 69 780 72
rect 744 63 747 69
rect 753 63 759 69
rect 765 63 771 69
rect 777 63 780 69
rect 744 60 780 63
rect 792 69 828 72
rect 792 63 795 69
rect 801 63 807 69
rect 813 63 819 69
rect 825 63 828 69
rect 792 60 828 63
rect 864 69 900 72
rect 864 63 867 69
rect 873 63 879 69
rect 885 63 891 69
rect 897 63 900 69
rect 864 60 900 63
rect 912 69 948 72
rect 912 63 915 69
rect 921 63 927 69
rect 933 63 939 69
rect 945 63 948 69
rect 912 60 948 63
rect 960 69 996 72
rect 960 63 963 69
rect 969 63 975 69
rect 981 63 987 69
rect 993 63 996 69
rect 960 60 996 63
rect 1008 69 1044 72
rect 1008 63 1011 69
rect 1017 63 1023 69
rect 1029 63 1035 69
rect 1041 63 1044 69
rect 1008 60 1044 63
rect 1080 69 1116 72
rect 1080 63 1083 69
rect 1089 63 1095 69
rect 1101 63 1107 69
rect 1113 63 1116 69
rect 1080 60 1116 63
rect 1128 69 1164 72
rect 1128 63 1131 69
rect 1137 63 1143 69
rect 1149 63 1155 69
rect 1161 63 1164 69
rect 1128 60 1164 63
rect 1176 69 1212 72
rect 1176 63 1179 69
rect 1185 63 1191 69
rect 1197 63 1203 69
rect 1209 63 1212 69
rect 1176 60 1212 63
rect 1224 69 1260 72
rect 1224 63 1227 69
rect 1233 63 1239 69
rect 1245 63 1251 69
rect 1257 63 1260 69
rect 1224 60 1260 63
rect 1296 69 1476 72
rect 1296 63 1299 69
rect 1305 63 1311 69
rect 1317 63 1323 69
rect 1329 63 1347 69
rect 1353 63 1359 69
rect 1365 63 1371 69
rect 1377 63 1395 69
rect 1401 63 1407 69
rect 1413 63 1419 69
rect 1425 63 1443 69
rect 1449 63 1455 69
rect 1461 63 1467 69
rect 1473 63 1476 69
rect 1296 60 1476 63
rect 1524 69 1536 75
rect 1524 63 1527 69
rect 1533 63 1536 69
rect -60 51 -57 57
rect -51 51 -48 57
rect -60 45 -48 51
rect -60 39 -57 45
rect -51 39 -48 45
rect -60 33 -48 39
rect -60 27 -57 33
rect -51 27 -48 33
rect -60 21 -48 27
rect -60 15 -57 21
rect -51 15 -48 21
rect -60 9 -48 15
rect -60 3 -57 9
rect -51 3 -48 9
rect -60 0 -48 3
rect -12 45 0 48
rect -12 39 -9 45
rect -3 39 0 45
rect -12 33 0 39
rect -12 27 -9 33
rect -3 27 0 33
rect -12 21 0 27
rect -12 15 -9 21
rect -3 15 0 21
rect -12 0 0 15
rect 36 45 48 48
rect 36 39 39 45
rect 45 39 48 45
rect 36 33 48 39
rect 36 27 39 33
rect 45 27 48 33
rect 36 21 48 27
rect 36 15 39 21
rect 45 15 48 21
rect 36 12 48 15
rect 84 45 96 48
rect 84 39 87 45
rect 93 39 96 45
rect 84 33 96 39
rect 84 27 87 33
rect 93 27 96 33
rect 84 21 96 27
rect 84 15 87 21
rect 93 15 96 21
rect 84 12 96 15
rect 132 45 144 48
rect 132 39 135 45
rect 141 39 144 45
rect 132 33 144 39
rect 132 27 135 33
rect 141 27 144 33
rect 132 21 144 27
rect 132 15 135 21
rect 141 15 144 21
rect 132 12 144 15
rect 180 45 192 48
rect 180 39 183 45
rect 189 39 192 45
rect 180 33 192 39
rect 180 27 183 33
rect 189 27 192 33
rect 180 21 192 27
rect 180 15 183 21
rect 189 15 192 21
rect 180 0 192 15
rect 204 45 216 48
rect 204 39 207 45
rect 213 39 216 45
rect 204 33 216 39
rect 204 27 207 33
rect 213 27 216 33
rect 204 21 216 27
rect 204 15 207 21
rect 213 15 216 21
rect 204 0 216 15
rect 252 45 264 48
rect 252 39 255 45
rect 261 39 264 45
rect 252 33 264 39
rect 252 27 255 33
rect 261 27 264 33
rect 252 21 264 27
rect 252 15 255 21
rect 261 15 264 21
rect 252 12 264 15
rect 300 45 312 48
rect 300 39 303 45
rect 309 39 312 45
rect 300 33 312 39
rect 300 27 303 33
rect 309 27 312 33
rect 300 21 312 27
rect 300 15 303 21
rect 309 15 312 21
rect 300 12 312 15
rect 348 45 360 48
rect 348 39 351 45
rect 357 39 360 45
rect 348 33 360 39
rect 348 27 351 33
rect 357 27 360 33
rect 348 21 360 27
rect 348 15 351 21
rect 357 15 360 21
rect 348 12 360 15
rect 396 45 408 48
rect 396 39 399 45
rect 405 39 408 45
rect 396 33 408 39
rect 396 27 399 33
rect 405 27 408 33
rect 396 21 408 27
rect 396 15 399 21
rect 405 15 408 21
rect 396 0 408 15
rect 420 45 432 48
rect 420 39 423 45
rect 429 39 432 45
rect 420 33 432 39
rect 420 27 423 33
rect 429 27 432 33
rect 420 21 432 27
rect 420 15 423 21
rect 429 15 432 21
rect 420 0 432 15
rect 516 45 528 48
rect 516 39 519 45
rect 525 39 528 45
rect 516 33 528 39
rect 516 27 519 33
rect 525 27 528 33
rect 516 21 528 27
rect 516 15 519 21
rect 525 15 528 21
rect 516 12 528 15
rect 612 45 624 48
rect 612 39 615 45
rect 621 39 624 45
rect 612 33 624 39
rect 612 27 615 33
rect 621 27 624 33
rect 612 21 624 27
rect 612 15 615 21
rect 621 15 624 21
rect 612 0 624 15
rect 636 45 648 48
rect 636 39 639 45
rect 645 39 648 45
rect 636 33 648 39
rect 636 27 639 33
rect 645 27 648 33
rect 636 21 648 27
rect 636 15 639 21
rect 645 15 648 21
rect 636 0 648 15
rect 732 45 744 48
rect 732 39 735 45
rect 741 39 744 45
rect 732 33 744 39
rect 732 27 735 33
rect 741 27 744 33
rect 732 21 744 27
rect 732 15 735 21
rect 741 15 744 21
rect 732 12 744 15
rect 828 45 840 48
rect 828 39 831 45
rect 837 39 840 45
rect 828 33 840 39
rect 828 27 831 33
rect 837 27 840 33
rect 828 21 840 27
rect 828 15 831 21
rect 837 15 840 21
rect 828 0 840 15
rect 852 45 864 48
rect 852 39 855 45
rect 861 39 864 45
rect 852 33 864 39
rect 852 27 855 33
rect 861 27 864 33
rect 852 21 864 27
rect 852 15 855 21
rect 861 15 864 21
rect 852 0 864 15
rect 1044 45 1056 48
rect 1044 39 1047 45
rect 1053 39 1056 45
rect 1044 33 1056 39
rect 1044 27 1047 33
rect 1053 27 1056 33
rect 1044 21 1056 27
rect 1044 15 1047 21
rect 1053 15 1056 21
rect 1044 12 1056 15
rect 1068 45 1080 48
rect 1068 39 1071 45
rect 1077 39 1080 45
rect 1068 33 1080 39
rect 1068 27 1071 33
rect 1077 27 1080 33
rect 1068 21 1080 27
rect 1068 15 1071 21
rect 1077 15 1080 21
rect 1068 0 1080 15
rect 1092 45 1104 48
rect 1092 39 1095 45
rect 1101 39 1104 45
rect 1092 33 1104 39
rect 1092 27 1095 33
rect 1101 27 1104 33
rect 1092 21 1104 27
rect 1092 15 1095 21
rect 1101 15 1104 21
rect 1092 12 1104 15
rect 1116 45 1128 48
rect 1116 39 1119 45
rect 1125 39 1128 45
rect 1116 33 1128 39
rect 1116 27 1119 33
rect 1125 27 1128 33
rect 1116 21 1128 27
rect 1116 15 1119 21
rect 1125 15 1128 21
rect 1116 0 1128 15
rect 1140 45 1152 48
rect 1140 39 1143 45
rect 1149 39 1152 45
rect 1140 33 1152 39
rect 1140 27 1143 33
rect 1149 27 1152 33
rect 1140 21 1152 27
rect 1140 15 1143 21
rect 1149 15 1152 21
rect 1140 12 1152 15
rect 1164 45 1176 48
rect 1164 39 1167 45
rect 1173 39 1176 45
rect 1164 33 1176 39
rect 1164 27 1167 33
rect 1173 27 1176 33
rect 1164 21 1176 27
rect 1164 15 1167 21
rect 1173 15 1176 21
rect 1164 0 1176 15
rect 1188 45 1200 48
rect 1188 39 1191 45
rect 1197 39 1200 45
rect 1188 33 1200 39
rect 1188 27 1191 33
rect 1197 27 1200 33
rect 1188 21 1200 27
rect 1188 15 1191 21
rect 1197 15 1200 21
rect 1188 12 1200 15
rect 1212 45 1224 48
rect 1212 39 1215 45
rect 1221 39 1224 45
rect 1212 33 1224 39
rect 1212 27 1215 33
rect 1221 27 1224 33
rect 1212 21 1224 27
rect 1212 15 1215 21
rect 1221 15 1224 21
rect 1212 0 1224 15
rect 1236 45 1248 48
rect 1236 39 1239 45
rect 1245 39 1248 45
rect 1236 33 1248 39
rect 1236 27 1239 33
rect 1245 27 1248 33
rect 1236 21 1248 27
rect 1236 15 1239 21
rect 1245 15 1248 21
rect 1236 12 1248 15
rect 1260 45 1272 48
rect 1260 39 1263 45
rect 1269 39 1272 45
rect 1260 33 1272 39
rect 1260 27 1263 33
rect 1269 27 1272 33
rect 1260 21 1272 27
rect 1260 15 1263 21
rect 1269 15 1272 21
rect 1260 0 1272 15
rect 1284 45 1296 48
rect 1284 39 1287 45
rect 1293 39 1296 45
rect 1284 33 1296 39
rect 1284 27 1287 33
rect 1293 27 1296 33
rect 1284 21 1296 27
rect 1284 15 1287 21
rect 1293 15 1296 21
rect 1284 0 1296 15
rect 1308 45 1320 60
rect 1308 39 1311 45
rect 1317 39 1320 45
rect 1308 33 1320 39
rect 1308 27 1311 33
rect 1317 27 1320 33
rect 1308 21 1320 27
rect 1308 15 1311 21
rect 1317 15 1320 21
rect 1308 12 1320 15
rect 1332 45 1344 48
rect 1332 39 1335 45
rect 1341 39 1344 45
rect 1332 33 1344 39
rect 1332 27 1335 33
rect 1341 27 1344 33
rect 1332 21 1344 27
rect 1332 15 1335 21
rect 1341 15 1344 21
rect 1332 0 1344 15
rect 1356 45 1368 60
rect 1356 39 1359 45
rect 1365 39 1368 45
rect 1356 33 1368 39
rect 1356 27 1359 33
rect 1365 27 1368 33
rect 1356 21 1368 27
rect 1356 15 1359 21
rect 1365 15 1368 21
rect 1356 12 1368 15
rect 1380 45 1392 48
rect 1380 39 1383 45
rect 1389 39 1392 45
rect 1380 33 1392 39
rect 1380 27 1383 33
rect 1389 27 1392 33
rect 1380 21 1392 27
rect 1380 15 1383 21
rect 1389 15 1392 21
rect 1380 0 1392 15
rect 1404 45 1416 60
rect 1404 39 1407 45
rect 1413 39 1416 45
rect 1404 33 1416 39
rect 1404 27 1407 33
rect 1413 27 1416 33
rect 1404 21 1416 27
rect 1404 15 1407 21
rect 1413 15 1416 21
rect 1404 12 1416 15
rect 1428 45 1440 48
rect 1428 39 1431 45
rect 1437 39 1440 45
rect 1428 33 1440 39
rect 1428 27 1431 33
rect 1437 27 1440 33
rect 1428 21 1440 27
rect 1428 15 1431 21
rect 1437 15 1440 21
rect 1428 0 1440 15
rect 1452 45 1464 60
rect 1524 57 1536 63
rect 1524 51 1527 57
rect 1533 51 1536 57
rect 1452 39 1455 45
rect 1461 39 1464 45
rect 1452 33 1464 39
rect 1452 27 1455 33
rect 1461 27 1464 33
rect 1452 21 1464 27
rect 1452 15 1455 21
rect 1461 15 1464 21
rect 1452 12 1464 15
rect 1476 45 1488 48
rect 1476 39 1479 45
rect 1485 39 1488 45
rect 1476 33 1488 39
rect 1476 27 1479 33
rect 1485 27 1488 33
rect 1476 21 1488 27
rect 1476 15 1479 21
rect 1485 15 1488 21
rect 1476 0 1488 15
rect 1524 45 1536 51
rect 1524 39 1527 45
rect 1533 39 1536 45
rect 1524 33 1536 39
rect 1524 27 1527 33
rect 1533 27 1536 33
rect 1524 21 1536 27
rect 1524 15 1527 21
rect 1533 15 1536 21
rect 1524 9 1536 15
rect 1524 3 1527 9
rect 1533 3 1536 9
rect 1524 0 1536 3
rect -60 -3 1536 0
rect -60 -9 -57 -3
rect -51 -9 -45 -3
rect -39 -9 -33 -3
rect -27 -9 -21 -3
rect -15 -9 -9 -3
rect -3 -9 3 -3
rect 9 -9 15 -3
rect 21 -9 27 -3
rect 33 -9 39 -3
rect 45 -9 51 -3
rect 57 -9 63 -3
rect 69 -9 75 -3
rect 81 -9 87 -3
rect 93 -9 99 -3
rect 105 -9 111 -3
rect 117 -9 123 -3
rect 129 -9 135 -3
rect 141 -9 147 -3
rect 153 -9 159 -3
rect 165 -9 171 -3
rect 177 -9 183 -3
rect 189 -9 195 -3
rect 201 -9 207 -3
rect 213 -9 219 -3
rect 225 -9 231 -3
rect 237 -9 243 -3
rect 249 -9 255 -3
rect 261 -9 267 -3
rect 273 -9 279 -3
rect 285 -9 291 -3
rect 297 -9 303 -3
rect 309 -9 315 -3
rect 321 -9 327 -3
rect 333 -9 339 -3
rect 345 -9 351 -3
rect 357 -9 363 -3
rect 369 -9 375 -3
rect 381 -9 387 -3
rect 393 -9 399 -3
rect 405 -9 411 -3
rect 417 -9 423 -3
rect 429 -9 435 -3
rect 441 -9 447 -3
rect 453 -9 459 -3
rect 465 -9 471 -3
rect 477 -9 483 -3
rect 489 -9 495 -3
rect 501 -9 507 -3
rect 513 -9 519 -3
rect 525 -9 531 -3
rect 537 -9 543 -3
rect 549 -9 555 -3
rect 561 -9 567 -3
rect 573 -9 579 -3
rect 585 -9 591 -3
rect 597 -9 603 -3
rect 609 -9 615 -3
rect 621 -9 627 -3
rect 633 -9 639 -3
rect 645 -9 651 -3
rect 657 -9 663 -3
rect 669 -9 675 -3
rect 681 -9 687 -3
rect 693 -9 699 -3
rect 705 -9 711 -3
rect 717 -9 723 -3
rect 729 -9 735 -3
rect 741 -9 747 -3
rect 753 -9 759 -3
rect 765 -9 771 -3
rect 777 -9 783 -3
rect 789 -9 795 -3
rect 801 -9 807 -3
rect 813 -9 819 -3
rect 825 -9 831 -3
rect 837 -9 843 -3
rect 849 -9 855 -3
rect 861 -9 867 -3
rect 873 -9 879 -3
rect 885 -9 891 -3
rect 897 -9 903 -3
rect 909 -9 915 -3
rect 921 -9 927 -3
rect 933 -9 939 -3
rect 945 -9 951 -3
rect 957 -9 963 -3
rect 969 -9 975 -3
rect 981 -9 987 -3
rect 993 -9 999 -3
rect 1005 -9 1011 -3
rect 1017 -9 1023 -3
rect 1029 -9 1035 -3
rect 1041 -9 1047 -3
rect 1053 -9 1059 -3
rect 1065 -9 1071 -3
rect 1077 -9 1083 -3
rect 1089 -9 1095 -3
rect 1101 -9 1107 -3
rect 1113 -9 1119 -3
rect 1125 -9 1131 -3
rect 1137 -9 1143 -3
rect 1149 -9 1155 -3
rect 1161 -9 1167 -3
rect 1173 -9 1179 -3
rect 1185 -9 1191 -3
rect 1197 -9 1203 -3
rect 1209 -9 1215 -3
rect 1221 -9 1227 -3
rect 1233 -9 1239 -3
rect 1245 -9 1251 -3
rect 1257 -9 1263 -3
rect 1269 -9 1275 -3
rect 1281 -9 1287 -3
rect 1293 -9 1299 -3
rect 1305 -9 1311 -3
rect 1317 -9 1323 -3
rect 1329 -9 1335 -3
rect 1341 -9 1347 -3
rect 1353 -9 1359 -3
rect 1365 -9 1371 -3
rect 1377 -9 1383 -3
rect 1389 -9 1395 -3
rect 1401 -9 1407 -3
rect 1413 -9 1419 -3
rect 1425 -9 1431 -3
rect 1437 -9 1443 -3
rect 1449 -9 1455 -3
rect 1461 -9 1467 -3
rect 1473 -9 1479 -3
rect 1485 -9 1491 -3
rect 1497 -9 1503 -3
rect 1509 -9 1515 -3
rect 1521 -9 1527 -3
rect 1533 -9 1536 -3
rect -60 -12 1536 -9
<< via1 >>
rect -9 567 -3 573
rect -9 555 -3 561
rect -9 543 -3 549
rect 15 567 21 573
rect 15 555 21 561
rect 15 543 21 549
rect 39 567 45 573
rect 39 555 45 561
rect 39 543 45 549
rect 63 567 69 573
rect 63 555 69 561
rect 63 543 69 549
rect 87 567 93 573
rect 87 555 93 561
rect 87 543 93 549
rect 111 567 117 573
rect 111 555 117 561
rect 111 543 117 549
rect 135 567 141 573
rect 135 555 141 561
rect 135 543 141 549
rect 159 567 165 573
rect 159 555 165 561
rect 159 543 165 549
rect 183 567 189 573
rect 183 555 189 561
rect 183 543 189 549
rect 207 567 213 573
rect 207 555 213 561
rect 207 543 213 549
rect 255 567 261 573
rect 255 555 261 561
rect 255 543 261 549
rect 303 567 309 573
rect 303 555 309 561
rect 303 543 309 549
rect 351 567 357 573
rect 351 555 357 561
rect 351 543 357 549
rect 399 567 405 573
rect 399 555 405 561
rect 399 543 405 549
rect 423 567 429 573
rect 423 555 429 561
rect 423 543 429 549
rect 471 567 477 573
rect 471 555 477 561
rect 471 543 477 549
rect 519 567 525 573
rect 519 555 525 561
rect 519 543 525 549
rect 567 567 573 573
rect 567 555 573 561
rect 567 543 573 549
rect 615 567 621 573
rect 615 555 621 561
rect 615 543 621 549
rect 639 567 645 573
rect 639 555 645 561
rect 639 543 645 549
rect 831 567 837 573
rect 831 555 837 561
rect 831 543 837 549
rect 855 567 861 573
rect 855 555 861 561
rect 855 543 861 549
rect 1047 567 1053 573
rect 1047 555 1053 561
rect 1047 543 1053 549
rect 1071 567 1077 573
rect 1071 555 1077 561
rect 1071 543 1077 549
rect 1095 567 1101 573
rect 1095 555 1101 561
rect 1095 543 1101 549
rect 1119 567 1125 573
rect 1119 555 1125 561
rect 1119 543 1125 549
rect 1143 567 1149 573
rect 1143 555 1149 561
rect 1143 543 1149 549
rect 1167 567 1173 573
rect 1167 555 1173 561
rect 1167 543 1173 549
rect 1191 567 1197 573
rect 1191 555 1197 561
rect 1191 543 1197 549
rect 1215 567 1221 573
rect 1215 555 1221 561
rect 1215 543 1221 549
rect 1239 567 1245 573
rect 1239 555 1245 561
rect 1239 543 1245 549
rect 1263 567 1269 573
rect 1263 555 1269 561
rect 1263 543 1269 549
rect 1287 567 1293 573
rect 1287 555 1293 561
rect 1287 543 1293 549
rect 1311 567 1317 573
rect 1311 555 1317 561
rect 1311 543 1317 549
rect 1335 567 1341 573
rect 1335 555 1341 561
rect 1335 543 1341 549
rect 1359 567 1365 573
rect 1359 555 1365 561
rect 1359 543 1365 549
rect 1383 567 1389 573
rect 1383 555 1389 561
rect 1383 543 1389 549
rect 1407 567 1413 573
rect 1407 555 1413 561
rect 1407 543 1413 549
rect 1431 567 1437 573
rect 1431 555 1437 561
rect 1431 543 1437 549
rect 1455 567 1461 573
rect 1455 555 1461 561
rect 1455 543 1461 549
rect 1479 567 1485 573
rect 1479 555 1485 561
rect 1479 543 1485 549
rect 39 519 45 525
rect 87 519 93 525
rect 135 519 141 525
rect 231 519 237 525
rect 279 519 285 525
rect 327 519 333 525
rect 375 519 381 525
rect 519 519 525 525
rect 639 519 645 525
rect 903 519 909 525
rect 1119 519 1125 525
rect 1167 519 1173 525
rect 1215 519 1221 525
rect 1335 519 1341 525
rect 1383 519 1389 525
rect 1431 519 1437 525
rect -9 471 -3 477
rect -9 459 -3 465
rect -9 447 -3 453
rect 15 471 21 477
rect 15 459 21 465
rect 15 447 21 453
rect 39 471 45 477
rect 39 459 45 465
rect 39 447 45 453
rect 63 471 69 477
rect 63 459 69 465
rect 63 447 69 453
rect 87 471 93 477
rect 87 459 93 465
rect 87 447 93 453
rect 111 471 117 477
rect 111 459 117 465
rect 111 447 117 453
rect 135 471 141 477
rect 135 459 141 465
rect 135 447 141 453
rect 159 471 165 477
rect 159 459 165 465
rect 159 447 165 453
rect 183 471 189 477
rect 183 459 189 465
rect 183 447 189 453
rect 207 471 213 477
rect 207 459 213 465
rect 207 447 213 453
rect 255 471 261 477
rect 255 459 261 465
rect 255 447 261 453
rect 303 471 309 477
rect 303 459 309 465
rect 303 447 309 453
rect 351 471 357 477
rect 351 459 357 465
rect 351 447 357 453
rect 399 471 405 477
rect 399 459 405 465
rect 399 447 405 453
rect 423 471 429 477
rect 423 459 429 465
rect 423 447 429 453
rect 471 471 477 477
rect 471 459 477 465
rect 471 447 477 453
rect 519 471 525 477
rect 519 459 525 465
rect 519 447 525 453
rect 567 471 573 477
rect 567 459 573 465
rect 567 447 573 453
rect 615 471 621 477
rect 615 459 621 465
rect 615 447 621 453
rect 639 471 645 477
rect 639 459 645 465
rect 639 447 645 453
rect 831 471 837 477
rect 831 459 837 465
rect 831 447 837 453
rect 855 471 861 477
rect 855 459 861 465
rect 855 447 861 453
rect 1047 471 1053 477
rect 1047 459 1053 465
rect 1047 447 1053 453
rect 1071 471 1077 477
rect 1071 459 1077 465
rect 1071 447 1077 453
rect 1095 471 1101 477
rect 1095 459 1101 465
rect 1095 447 1101 453
rect 1119 471 1125 477
rect 1119 459 1125 465
rect 1119 447 1125 453
rect 1143 471 1149 477
rect 1143 459 1149 465
rect 1143 447 1149 453
rect 1167 471 1173 477
rect 1167 459 1173 465
rect 1167 447 1173 453
rect 1191 471 1197 477
rect 1191 459 1197 465
rect 1191 447 1197 453
rect 1215 471 1221 477
rect 1215 459 1221 465
rect 1215 447 1221 453
rect 1239 471 1245 477
rect 1239 459 1245 465
rect 1239 447 1245 453
rect 1263 471 1269 477
rect 1263 459 1269 465
rect 1263 447 1269 453
rect 1287 471 1293 477
rect 1287 459 1293 465
rect 1287 447 1293 453
rect 1311 471 1317 477
rect 1311 459 1317 465
rect 1311 447 1317 453
rect 1335 471 1341 477
rect 1335 459 1341 465
rect 1335 447 1341 453
rect 1359 471 1365 477
rect 1359 459 1365 465
rect 1359 447 1365 453
rect 1383 471 1389 477
rect 1383 459 1389 465
rect 1383 447 1389 453
rect 1407 471 1413 477
rect 1407 459 1413 465
rect 1407 447 1413 453
rect 1431 471 1437 477
rect 1431 459 1437 465
rect 1431 447 1437 453
rect 1455 471 1461 477
rect 1455 459 1461 465
rect 1455 447 1461 453
rect 1479 471 1485 477
rect 1479 459 1485 465
rect 1479 447 1485 453
rect 15 423 21 429
rect 63 423 69 429
rect 111 423 117 429
rect 159 423 165 429
rect 231 423 237 429
rect 279 423 285 429
rect 327 423 333 429
rect 375 423 381 429
rect 447 423 453 429
rect 495 423 501 429
rect 543 423 549 429
rect 591 423 597 429
rect 639 423 645 429
rect 663 423 669 429
rect 711 423 717 429
rect 759 423 765 429
rect 807 423 813 429
rect 831 423 837 429
rect 903 423 909 429
rect 1095 423 1101 429
rect 1143 423 1149 429
rect 1191 423 1197 429
rect 1239 423 1245 429
rect 1311 423 1317 429
rect 1359 423 1365 429
rect 1407 423 1413 429
rect 1455 423 1461 429
rect -33 399 -27 405
rect -33 351 -27 357
rect -9 303 -3 309
rect 39 303 45 309
rect 87 303 93 309
rect 135 303 141 309
rect 183 303 189 309
rect 231 303 237 309
rect 279 303 285 309
rect 327 303 333 309
rect 375 303 381 309
rect 447 303 453 309
rect 495 303 501 309
rect 543 303 549 309
rect 591 303 597 309
rect 663 303 669 309
rect 711 303 717 309
rect 759 303 765 309
rect 807 303 813 309
rect 867 303 873 309
rect 927 303 933 309
rect 975 303 981 309
rect 1023 303 1029 309
rect 1095 303 1101 309
rect 1143 303 1149 309
rect 1191 303 1197 309
rect 1239 303 1245 309
rect 1311 303 1317 309
rect 1359 303 1365 309
rect 1407 303 1413 309
rect 1455 303 1461 309
rect -9 279 -3 285
rect -9 267 -3 273
rect -9 255 -3 261
rect 39 279 45 285
rect 39 267 45 273
rect 39 255 45 261
rect 87 279 93 285
rect 87 267 93 273
rect 87 255 93 261
rect 135 279 141 285
rect 135 267 141 273
rect 135 255 141 261
rect 183 279 189 285
rect 183 267 189 273
rect 183 255 189 261
rect 207 279 213 285
rect 207 267 213 273
rect 207 255 213 261
rect 303 279 309 285
rect 303 267 309 273
rect 303 255 309 261
rect 399 279 405 285
rect 399 267 405 273
rect 399 255 405 261
rect 423 279 429 285
rect 423 267 429 273
rect 423 255 429 261
rect 519 279 525 285
rect 519 267 525 273
rect 519 255 525 261
rect 615 279 621 285
rect 615 267 621 273
rect 615 255 621 261
rect 639 279 645 285
rect 639 267 645 273
rect 639 255 645 261
rect 735 279 741 285
rect 735 267 741 273
rect 735 255 741 261
rect 831 279 837 285
rect 831 267 837 273
rect 831 255 837 261
rect 855 279 861 285
rect 855 267 861 273
rect 855 255 861 261
rect 879 279 885 285
rect 879 267 885 273
rect 879 255 885 261
rect 903 279 909 285
rect 903 267 909 273
rect 903 255 909 261
rect 1047 279 1053 285
rect 1047 267 1053 273
rect 1047 255 1053 261
rect 1071 279 1077 285
rect 1071 267 1077 273
rect 1071 255 1077 261
rect 1095 255 1101 261
rect 1119 279 1125 285
rect 1143 255 1149 261
rect 1167 279 1173 285
rect 1191 255 1197 261
rect 1215 279 1221 285
rect 1239 255 1245 261
rect 1263 279 1269 285
rect 1263 267 1269 273
rect 1263 255 1269 261
rect 1287 279 1293 285
rect 1287 267 1293 273
rect 1287 255 1293 261
rect 1311 255 1317 261
rect 1335 279 1341 285
rect 1359 255 1365 261
rect 1383 279 1389 285
rect 1407 255 1413 261
rect 1431 279 1437 285
rect 1455 255 1461 261
rect 1479 279 1485 285
rect 1479 267 1485 273
rect 1479 255 1485 261
rect -57 207 -51 213
rect 1527 207 1533 213
rect 15 63 21 69
rect 63 63 69 69
rect 111 63 117 69
rect 159 63 165 69
rect 231 63 237 69
rect 279 63 285 69
rect 327 63 333 69
rect 375 63 381 69
rect 447 63 453 69
rect 495 63 501 69
rect 543 63 549 69
rect 591 63 597 69
rect 663 63 669 69
rect 711 63 717 69
rect 759 63 765 69
rect 807 63 813 69
rect 879 63 885 69
rect 927 63 933 69
rect 975 63 981 69
rect 1023 63 1029 69
rect 1095 63 1101 69
rect 1143 63 1149 69
rect 1191 63 1197 69
rect 1239 63 1245 69
rect -9 39 -3 45
rect -9 27 -3 33
rect -9 15 -3 21
rect 39 39 45 45
rect 39 27 45 33
rect 39 15 45 21
rect 87 39 93 45
rect 87 27 93 33
rect 87 15 93 21
rect 135 39 141 45
rect 135 27 141 33
rect 135 15 141 21
rect 183 39 189 45
rect 183 27 189 33
rect 183 15 189 21
rect 207 39 213 45
rect 207 27 213 33
rect 207 15 213 21
rect 255 39 261 45
rect 255 27 261 33
rect 255 15 261 21
rect 303 39 309 45
rect 303 27 309 33
rect 303 15 309 21
rect 351 39 357 45
rect 351 27 357 33
rect 351 15 357 21
rect 399 39 405 45
rect 399 27 405 33
rect 399 15 405 21
rect 423 39 429 45
rect 423 27 429 33
rect 423 15 429 21
rect 519 39 525 45
rect 519 27 525 33
rect 519 15 525 21
rect 615 39 621 45
rect 615 27 621 33
rect 615 15 621 21
rect 639 39 645 45
rect 639 27 645 33
rect 639 15 645 21
rect 735 39 741 45
rect 735 27 741 33
rect 735 15 741 21
rect 831 39 837 45
rect 831 27 837 33
rect 831 15 837 21
rect 855 39 861 45
rect 855 27 861 33
rect 855 15 861 21
rect 1047 39 1053 45
rect 1047 27 1053 33
rect 1047 15 1053 21
rect 1071 39 1077 45
rect 1071 27 1077 33
rect 1071 15 1077 21
rect 1095 39 1101 45
rect 1119 15 1125 21
rect 1143 39 1149 45
rect 1167 39 1173 45
rect 1167 27 1173 33
rect 1167 15 1173 21
rect 1191 39 1197 45
rect 1215 15 1221 21
rect 1239 39 1245 45
rect 1263 39 1269 45
rect 1263 27 1269 33
rect 1263 15 1269 21
<< metal2 >>
rect -12 573 0 576
rect -12 567 -9 573
rect -3 567 0 573
rect -12 561 0 567
rect -12 555 -9 561
rect -3 555 0 561
rect -12 549 0 555
rect -12 543 -9 549
rect -3 543 0 549
rect -12 501 0 543
rect -12 495 -9 501
rect -3 495 0 501
rect -12 492 0 495
rect 12 573 24 576
rect 12 567 15 573
rect 21 567 24 573
rect 12 561 24 567
rect 12 555 15 561
rect 21 555 24 561
rect 12 549 24 555
rect 12 543 15 549
rect 21 543 24 549
rect -12 477 0 480
rect -12 471 -9 477
rect -3 471 0 477
rect -12 465 0 471
rect -12 459 -9 465
rect -3 459 0 465
rect -12 453 0 459
rect -12 447 -9 453
rect -3 447 0 453
rect -36 405 -24 408
rect -36 399 -33 405
rect -27 399 -24 405
rect -36 396 -24 399
rect -36 357 -24 360
rect -36 351 -33 357
rect -27 351 -24 357
rect -36 348 -24 351
rect -12 309 0 447
rect 12 477 24 543
rect 36 573 48 576
rect 36 567 39 573
rect 45 567 48 573
rect 36 561 48 567
rect 36 555 39 561
rect 45 555 48 561
rect 36 549 48 555
rect 36 543 39 549
rect 45 543 48 549
rect 36 540 48 543
rect 60 573 72 576
rect 60 567 63 573
rect 69 567 72 573
rect 60 561 72 567
rect 60 555 63 561
rect 69 555 72 561
rect 60 549 72 555
rect 60 543 63 549
rect 69 543 72 549
rect 36 525 48 528
rect 36 519 39 525
rect 45 519 48 525
rect 36 516 48 519
rect 12 471 15 477
rect 21 471 24 477
rect 12 465 24 471
rect 12 459 15 465
rect 21 459 24 465
rect 12 453 24 459
rect 12 447 15 453
rect 21 447 24 453
rect 12 444 24 447
rect 36 477 48 480
rect 36 471 39 477
rect 45 471 48 477
rect 36 465 48 471
rect 36 459 39 465
rect 45 459 48 465
rect 36 453 48 459
rect 36 447 39 453
rect 45 447 48 453
rect 12 429 24 432
rect 12 423 15 429
rect 21 423 24 429
rect 12 420 24 423
rect -12 303 -9 309
rect -3 303 0 309
rect -12 300 0 303
rect 12 300 24 312
rect 36 309 48 447
rect 60 477 72 543
rect 84 573 96 576
rect 84 567 87 573
rect 93 567 96 573
rect 84 561 96 567
rect 84 555 87 561
rect 93 555 96 561
rect 84 549 96 555
rect 84 543 87 549
rect 93 543 96 549
rect 84 540 96 543
rect 108 573 120 576
rect 108 567 111 573
rect 117 567 120 573
rect 108 561 120 567
rect 108 555 111 561
rect 117 555 120 561
rect 108 549 120 555
rect 108 543 111 549
rect 117 543 120 549
rect 84 525 96 528
rect 84 519 87 525
rect 93 519 96 525
rect 84 516 96 519
rect 60 471 63 477
rect 69 471 72 477
rect 60 465 72 471
rect 60 459 63 465
rect 69 459 72 465
rect 60 453 72 459
rect 60 447 63 453
rect 69 447 72 453
rect 60 444 72 447
rect 84 477 96 480
rect 84 471 87 477
rect 93 471 96 477
rect 84 465 96 471
rect 84 459 87 465
rect 93 459 96 465
rect 84 453 96 459
rect 84 447 87 453
rect 93 447 96 453
rect 60 429 72 432
rect 60 423 63 429
rect 69 423 72 429
rect 60 420 72 423
rect 36 303 39 309
rect 45 303 48 309
rect 36 300 48 303
rect 60 300 72 312
rect 84 309 96 447
rect 108 477 120 543
rect 132 573 144 576
rect 132 567 135 573
rect 141 567 144 573
rect 132 561 144 567
rect 132 555 135 561
rect 141 555 144 561
rect 132 549 144 555
rect 132 543 135 549
rect 141 543 144 549
rect 132 540 144 543
rect 156 573 168 576
rect 156 567 159 573
rect 165 567 168 573
rect 156 561 168 567
rect 156 555 159 561
rect 165 555 168 561
rect 156 549 168 555
rect 156 543 159 549
rect 165 543 168 549
rect 132 525 144 528
rect 132 519 135 525
rect 141 519 144 525
rect 132 516 144 519
rect 108 471 111 477
rect 117 471 120 477
rect 108 465 120 471
rect 108 459 111 465
rect 117 459 120 465
rect 108 453 120 459
rect 108 447 111 453
rect 117 447 120 453
rect 108 444 120 447
rect 132 477 144 480
rect 132 471 135 477
rect 141 471 144 477
rect 132 465 144 471
rect 132 459 135 465
rect 141 459 144 465
rect 132 453 144 459
rect 132 447 135 453
rect 141 447 144 453
rect 108 429 120 432
rect 108 423 111 429
rect 117 423 120 429
rect 108 420 120 423
rect 84 303 87 309
rect 93 303 96 309
rect 84 300 96 303
rect 132 309 144 447
rect 156 477 168 543
rect 180 573 192 576
rect 180 567 183 573
rect 189 567 192 573
rect 180 561 192 567
rect 180 555 183 561
rect 189 555 192 561
rect 180 549 192 555
rect 180 543 183 549
rect 189 543 192 549
rect 180 540 192 543
rect 204 573 216 576
rect 204 567 207 573
rect 213 567 216 573
rect 204 561 216 567
rect 204 555 207 561
rect 213 555 216 561
rect 204 549 216 555
rect 204 543 207 549
rect 213 543 216 549
rect 204 540 216 543
rect 252 573 264 576
rect 252 567 255 573
rect 261 567 264 573
rect 252 561 264 567
rect 252 555 255 561
rect 261 555 264 561
rect 252 549 264 555
rect 252 543 255 549
rect 261 543 264 549
rect 228 525 240 528
rect 228 519 231 525
rect 237 519 240 525
rect 228 516 240 519
rect 156 471 159 477
rect 165 471 168 477
rect 156 465 168 471
rect 156 459 159 465
rect 165 459 168 465
rect 156 453 168 459
rect 156 447 159 453
rect 165 447 168 453
rect 156 444 168 447
rect 180 477 192 480
rect 180 471 183 477
rect 189 471 192 477
rect 180 465 192 471
rect 180 459 183 465
rect 189 459 192 465
rect 180 453 192 459
rect 180 447 183 453
rect 189 447 192 453
rect 156 429 168 432
rect 156 423 159 429
rect 165 423 168 429
rect 156 420 168 423
rect 132 303 135 309
rect 141 303 144 309
rect 132 300 144 303
rect 180 309 192 447
rect 180 303 183 309
rect 189 303 192 309
rect 180 300 192 303
rect 204 477 216 480
rect 204 471 207 477
rect 213 471 216 477
rect 204 465 216 471
rect 204 459 207 465
rect 213 459 216 465
rect 204 453 216 459
rect 204 447 207 453
rect 213 447 216 453
rect -12 285 0 288
rect -12 279 -9 285
rect -3 279 0 285
rect -12 273 0 279
rect -12 267 -9 273
rect -3 267 0 273
rect -12 261 0 267
rect -12 255 -9 261
rect -3 255 0 261
rect -60 213 -48 216
rect -60 207 -57 213
rect -51 207 -48 213
rect -60 204 -48 207
rect -12 189 0 255
rect -12 183 -9 189
rect -3 183 0 189
rect -12 180 0 183
rect 36 285 48 288
rect 36 279 39 285
rect 45 279 48 285
rect 36 273 48 279
rect 36 267 39 273
rect 45 267 48 273
rect 36 261 48 267
rect 36 255 39 261
rect 45 255 48 261
rect 36 189 48 255
rect 36 183 39 189
rect 45 183 48 189
rect 36 180 48 183
rect 84 285 96 288
rect 84 279 87 285
rect 93 279 96 285
rect 84 273 96 279
rect 84 267 87 273
rect 93 267 96 273
rect 84 261 96 267
rect 84 255 87 261
rect 93 255 96 261
rect 84 189 96 255
rect 84 183 87 189
rect 93 183 96 189
rect 36 165 48 168
rect 36 159 39 165
rect 45 159 48 165
rect 12 69 24 72
rect 12 63 15 69
rect 21 63 24 69
rect 12 60 24 63
rect -12 45 0 48
rect -12 39 -9 45
rect -3 39 0 45
rect -12 33 0 39
rect -12 27 -9 33
rect -3 27 0 33
rect -12 21 0 27
rect -12 15 -9 21
rect -3 15 0 21
rect -12 12 0 15
rect 36 45 48 159
rect 60 69 72 72
rect 60 63 63 69
rect 69 63 72 69
rect 60 60 72 63
rect 36 39 39 45
rect 45 39 48 45
rect 36 33 48 39
rect 36 27 39 33
rect 45 27 48 33
rect 36 21 48 27
rect 36 15 39 21
rect 45 15 48 21
rect 36 12 48 15
rect 84 45 96 183
rect 132 285 144 288
rect 132 279 135 285
rect 141 279 144 285
rect 132 273 144 279
rect 132 267 135 273
rect 141 267 144 273
rect 132 261 144 267
rect 132 255 135 261
rect 141 255 144 261
rect 132 189 144 255
rect 132 183 135 189
rect 141 183 144 189
rect 132 180 144 183
rect 180 285 192 288
rect 180 279 183 285
rect 189 279 192 285
rect 180 273 192 279
rect 180 267 183 273
rect 189 267 192 273
rect 180 261 192 267
rect 180 255 183 261
rect 189 255 192 261
rect 180 189 192 255
rect 204 285 216 447
rect 252 477 264 543
rect 300 573 312 576
rect 300 567 303 573
rect 309 567 312 573
rect 300 561 312 567
rect 300 555 303 561
rect 309 555 312 561
rect 300 549 312 555
rect 300 543 303 549
rect 309 543 312 549
rect 300 540 312 543
rect 348 573 360 576
rect 348 567 351 573
rect 357 567 360 573
rect 348 561 360 567
rect 348 555 351 561
rect 357 555 360 561
rect 348 549 360 555
rect 348 543 351 549
rect 357 543 360 549
rect 276 525 288 528
rect 276 519 279 525
rect 285 519 288 525
rect 276 516 288 519
rect 324 525 336 528
rect 324 519 327 525
rect 333 519 336 525
rect 324 516 336 519
rect 252 471 255 477
rect 261 471 264 477
rect 252 465 264 471
rect 252 459 255 465
rect 261 459 264 465
rect 252 453 264 459
rect 252 447 255 453
rect 261 447 264 453
rect 252 444 264 447
rect 300 477 312 480
rect 300 471 303 477
rect 309 471 312 477
rect 300 465 312 471
rect 300 459 303 465
rect 309 459 312 465
rect 300 453 312 459
rect 300 447 303 453
rect 309 447 312 453
rect 300 444 312 447
rect 348 477 360 543
rect 396 573 408 576
rect 396 567 399 573
rect 405 567 408 573
rect 396 561 408 567
rect 396 555 399 561
rect 405 555 408 561
rect 396 549 408 555
rect 396 543 399 549
rect 405 543 408 549
rect 396 540 408 543
rect 420 573 432 576
rect 420 567 423 573
rect 429 567 432 573
rect 420 561 432 567
rect 420 555 423 561
rect 429 555 432 561
rect 420 549 432 555
rect 420 543 423 549
rect 429 543 432 549
rect 420 540 432 543
rect 468 573 480 576
rect 468 567 471 573
rect 477 567 480 573
rect 468 561 480 567
rect 468 555 471 561
rect 477 555 480 561
rect 468 549 480 555
rect 468 543 471 549
rect 477 543 480 549
rect 372 525 384 528
rect 372 519 375 525
rect 381 519 384 525
rect 372 516 384 519
rect 348 471 351 477
rect 357 471 360 477
rect 348 465 360 471
rect 348 459 351 465
rect 357 459 360 465
rect 348 453 360 459
rect 348 447 351 453
rect 357 447 360 453
rect 348 444 360 447
rect 396 477 408 480
rect 396 471 399 477
rect 405 471 408 477
rect 396 465 408 471
rect 396 459 399 465
rect 405 459 408 465
rect 396 453 408 459
rect 396 447 399 453
rect 405 447 408 453
rect 228 429 240 432
rect 228 423 231 429
rect 237 423 240 429
rect 228 420 240 423
rect 276 429 288 432
rect 276 423 279 429
rect 285 423 288 429
rect 276 420 288 423
rect 324 429 336 432
rect 324 423 327 429
rect 333 423 336 429
rect 324 420 336 423
rect 372 429 384 432
rect 372 423 375 429
rect 381 423 384 429
rect 372 420 384 423
rect 228 309 240 312
rect 228 303 231 309
rect 237 303 240 309
rect 228 300 240 303
rect 276 309 288 312
rect 276 303 279 309
rect 285 303 288 309
rect 276 300 288 303
rect 324 309 336 312
rect 324 303 327 309
rect 333 303 336 309
rect 324 300 336 303
rect 372 309 384 312
rect 372 303 375 309
rect 381 303 384 309
rect 372 300 384 303
rect 204 279 207 285
rect 213 279 216 285
rect 204 273 216 279
rect 204 267 207 273
rect 213 267 216 273
rect 204 261 216 267
rect 204 255 207 261
rect 213 255 216 261
rect 204 252 216 255
rect 300 285 312 288
rect 300 279 303 285
rect 309 279 312 285
rect 300 273 312 279
rect 300 267 303 273
rect 309 267 312 273
rect 300 261 312 267
rect 300 255 303 261
rect 309 255 312 261
rect 252 204 264 216
rect 180 183 183 189
rect 189 183 192 189
rect 180 180 192 183
rect 132 165 144 168
rect 132 159 135 165
rect 141 159 144 165
rect 108 69 120 72
rect 108 63 111 69
rect 117 63 120 69
rect 108 60 120 63
rect 84 39 87 45
rect 93 39 96 45
rect 84 33 96 39
rect 84 27 87 33
rect 93 27 96 33
rect 84 21 96 27
rect 84 15 87 21
rect 93 15 96 21
rect 84 12 96 15
rect 132 45 144 159
rect 252 165 264 168
rect 252 159 255 165
rect 261 159 264 165
rect 156 69 168 72
rect 156 63 159 69
rect 165 63 168 69
rect 156 60 168 63
rect 228 69 240 72
rect 228 63 231 69
rect 237 63 240 69
rect 228 60 240 63
rect 132 39 135 45
rect 141 39 144 45
rect 132 33 144 39
rect 132 27 135 33
rect 141 27 144 33
rect 132 21 144 27
rect 132 15 135 21
rect 141 15 144 21
rect 132 12 144 15
rect 180 45 192 48
rect 180 39 183 45
rect 189 39 192 45
rect 180 33 192 39
rect 180 27 183 33
rect 189 27 192 33
rect 180 21 192 27
rect 180 15 183 21
rect 189 15 192 21
rect 180 12 192 15
rect 204 45 216 48
rect 204 39 207 45
rect 213 39 216 45
rect 204 33 216 39
rect 204 27 207 33
rect 213 27 216 33
rect 204 21 216 27
rect 204 15 207 21
rect 213 15 216 21
rect 204 12 216 15
rect 252 45 264 159
rect 300 141 312 255
rect 396 285 408 447
rect 396 279 399 285
rect 405 279 408 285
rect 396 273 408 279
rect 396 267 399 273
rect 405 267 408 273
rect 396 261 408 267
rect 396 255 399 261
rect 405 255 408 261
rect 396 252 408 255
rect 420 477 432 480
rect 420 471 423 477
rect 429 471 432 477
rect 420 465 432 471
rect 420 459 423 465
rect 429 459 432 465
rect 420 453 432 459
rect 420 447 423 453
rect 429 447 432 453
rect 420 309 432 447
rect 468 477 480 543
rect 516 573 528 576
rect 516 567 519 573
rect 525 567 528 573
rect 516 561 528 567
rect 516 555 519 561
rect 525 555 528 561
rect 516 549 528 555
rect 516 543 519 549
rect 525 543 528 549
rect 516 540 528 543
rect 564 573 576 576
rect 564 567 567 573
rect 573 567 576 573
rect 564 561 576 567
rect 564 555 567 561
rect 573 555 576 561
rect 564 549 576 555
rect 564 543 567 549
rect 573 543 576 549
rect 516 525 528 528
rect 516 519 519 525
rect 525 519 528 525
rect 516 516 528 519
rect 468 471 471 477
rect 477 471 480 477
rect 468 465 480 471
rect 468 459 471 465
rect 477 459 480 465
rect 468 453 480 459
rect 468 447 471 453
rect 477 447 480 453
rect 468 444 480 447
rect 516 477 528 480
rect 516 471 519 477
rect 525 471 528 477
rect 516 465 528 471
rect 516 459 519 465
rect 525 459 528 465
rect 516 453 528 459
rect 516 447 519 453
rect 525 447 528 453
rect 516 444 528 447
rect 564 477 576 543
rect 612 573 624 576
rect 612 567 615 573
rect 621 567 624 573
rect 612 561 624 567
rect 612 555 615 561
rect 621 555 624 561
rect 612 549 624 555
rect 612 543 615 549
rect 621 543 624 549
rect 612 540 624 543
rect 636 573 648 576
rect 636 567 639 573
rect 645 567 648 573
rect 636 561 648 567
rect 636 555 639 561
rect 645 555 648 561
rect 636 549 648 555
rect 636 543 639 549
rect 645 543 648 549
rect 636 540 648 543
rect 828 573 840 576
rect 828 567 831 573
rect 837 567 840 573
rect 828 561 840 567
rect 828 555 831 561
rect 837 555 840 561
rect 828 549 840 555
rect 828 543 831 549
rect 837 543 840 549
rect 636 525 648 528
rect 636 519 639 525
rect 645 519 648 525
rect 564 471 567 477
rect 573 471 576 477
rect 564 465 576 471
rect 564 459 567 465
rect 573 459 576 465
rect 564 453 576 459
rect 564 447 567 453
rect 573 447 576 453
rect 564 444 576 447
rect 612 477 624 480
rect 612 471 615 477
rect 621 471 624 477
rect 612 465 624 471
rect 612 459 615 465
rect 621 459 624 465
rect 612 453 624 459
rect 612 447 615 453
rect 621 447 624 453
rect 444 429 456 432
rect 444 423 447 429
rect 453 423 456 429
rect 444 420 456 423
rect 492 429 504 432
rect 492 423 495 429
rect 501 423 504 429
rect 492 420 504 423
rect 540 429 552 432
rect 540 423 543 429
rect 549 423 552 429
rect 540 420 552 423
rect 588 429 600 432
rect 588 423 591 429
rect 597 423 600 429
rect 588 420 600 423
rect 420 303 423 309
rect 429 303 432 309
rect 420 285 432 303
rect 444 309 456 312
rect 444 303 447 309
rect 453 303 456 309
rect 444 300 456 303
rect 492 309 504 312
rect 492 303 495 309
rect 501 303 504 309
rect 492 300 504 303
rect 540 309 552 312
rect 540 303 543 309
rect 549 303 552 309
rect 540 300 552 303
rect 588 309 600 312
rect 588 303 591 309
rect 597 303 600 309
rect 588 300 600 303
rect 420 279 423 285
rect 429 279 432 285
rect 420 273 432 279
rect 420 267 423 273
rect 429 267 432 273
rect 420 261 432 267
rect 420 255 423 261
rect 429 255 432 261
rect 420 252 432 255
rect 516 285 528 288
rect 516 279 519 285
rect 525 279 528 285
rect 516 273 528 279
rect 516 267 519 273
rect 525 267 528 273
rect 516 261 528 267
rect 516 255 519 261
rect 525 255 528 261
rect 348 204 360 216
rect 300 135 303 141
rect 309 135 312 141
rect 276 69 288 72
rect 276 63 279 69
rect 285 63 288 69
rect 276 60 288 63
rect 252 39 255 45
rect 261 39 264 45
rect 252 33 264 39
rect 252 27 255 33
rect 261 27 264 33
rect 252 21 264 27
rect 252 15 255 21
rect 261 15 264 21
rect 252 12 264 15
rect 300 45 312 135
rect 348 165 360 168
rect 348 159 351 165
rect 357 159 360 165
rect 324 69 336 72
rect 324 63 327 69
rect 333 63 336 69
rect 324 60 336 63
rect 300 39 303 45
rect 309 39 312 45
rect 300 33 312 39
rect 300 27 303 33
rect 309 27 312 33
rect 300 21 312 27
rect 300 15 303 21
rect 309 15 312 21
rect 300 12 312 15
rect 348 45 360 159
rect 516 117 528 255
rect 612 285 624 447
rect 612 279 615 285
rect 621 279 624 285
rect 612 273 624 279
rect 612 267 615 273
rect 621 267 624 273
rect 612 261 624 267
rect 612 255 615 261
rect 621 255 624 261
rect 612 252 624 255
rect 636 477 648 519
rect 636 471 639 477
rect 645 471 648 477
rect 636 465 648 471
rect 636 459 639 465
rect 645 459 648 465
rect 636 453 648 459
rect 636 447 639 453
rect 645 447 648 453
rect 636 429 648 447
rect 828 477 840 543
rect 828 471 831 477
rect 837 471 840 477
rect 828 465 840 471
rect 828 459 831 465
rect 837 459 840 465
rect 828 453 840 459
rect 828 447 831 453
rect 837 447 840 453
rect 828 444 840 447
rect 852 573 864 576
rect 852 567 855 573
rect 861 567 864 573
rect 852 561 864 567
rect 852 555 855 561
rect 861 555 864 561
rect 852 549 864 555
rect 852 543 855 549
rect 861 543 864 549
rect 852 477 864 543
rect 1044 573 1056 576
rect 1044 567 1047 573
rect 1053 567 1056 573
rect 1044 561 1056 567
rect 1044 555 1047 561
rect 1053 555 1056 561
rect 1044 549 1056 555
rect 1044 543 1047 549
rect 1053 543 1056 549
rect 852 471 855 477
rect 861 471 864 477
rect 852 465 864 471
rect 852 459 855 465
rect 861 459 864 465
rect 852 453 864 459
rect 852 447 855 453
rect 861 447 864 453
rect 852 444 864 447
rect 900 525 912 528
rect 900 519 903 525
rect 909 519 912 525
rect 636 423 639 429
rect 645 423 648 429
rect 636 285 648 423
rect 660 429 672 432
rect 660 423 663 429
rect 669 423 672 429
rect 660 420 672 423
rect 708 429 720 432
rect 708 423 711 429
rect 717 423 720 429
rect 708 420 720 423
rect 756 429 768 432
rect 756 423 759 429
rect 765 423 768 429
rect 756 420 768 423
rect 804 429 816 432
rect 804 423 807 429
rect 813 423 816 429
rect 804 420 816 423
rect 828 429 840 432
rect 828 423 831 429
rect 837 423 840 429
rect 660 309 672 312
rect 660 303 663 309
rect 669 303 672 309
rect 660 300 672 303
rect 708 309 720 312
rect 708 303 711 309
rect 717 303 720 309
rect 708 300 720 303
rect 756 309 768 312
rect 756 303 759 309
rect 765 303 768 309
rect 756 300 768 303
rect 804 309 816 312
rect 804 303 807 309
rect 813 303 816 309
rect 804 300 816 303
rect 636 279 639 285
rect 645 279 648 285
rect 636 273 648 279
rect 636 267 639 273
rect 645 267 648 273
rect 636 261 648 267
rect 636 255 639 261
rect 645 255 648 261
rect 636 252 648 255
rect 732 285 744 288
rect 732 279 735 285
rect 741 279 744 285
rect 732 273 744 279
rect 732 267 735 273
rect 741 267 744 273
rect 732 261 744 267
rect 732 255 735 261
rect 741 255 744 261
rect 516 111 519 117
rect 525 111 528 117
rect 372 69 384 72
rect 372 63 375 69
rect 381 63 384 69
rect 372 60 384 63
rect 444 69 456 72
rect 444 63 447 69
rect 453 63 456 69
rect 444 60 456 63
rect 492 69 504 72
rect 492 63 495 69
rect 501 63 504 69
rect 492 60 504 63
rect 348 39 351 45
rect 357 39 360 45
rect 348 33 360 39
rect 348 27 351 33
rect 357 27 360 33
rect 348 21 360 27
rect 348 15 351 21
rect 357 15 360 21
rect 348 12 360 15
rect 396 45 408 48
rect 396 39 399 45
rect 405 39 408 45
rect 396 33 408 39
rect 396 27 399 33
rect 405 27 408 33
rect 396 21 408 27
rect 396 15 399 21
rect 405 15 408 21
rect 396 12 408 15
rect 420 45 432 48
rect 420 39 423 45
rect 429 39 432 45
rect 420 33 432 39
rect 420 27 423 33
rect 429 27 432 33
rect 420 21 432 27
rect 420 15 423 21
rect 429 15 432 21
rect 420 12 432 15
rect 516 45 528 111
rect 540 69 552 72
rect 540 63 543 69
rect 549 63 552 69
rect 540 60 552 63
rect 588 69 600 72
rect 588 63 591 69
rect 597 63 600 69
rect 588 60 600 63
rect 660 69 672 72
rect 660 63 663 69
rect 669 63 672 69
rect 660 60 672 63
rect 708 69 720 72
rect 708 63 711 69
rect 717 63 720 69
rect 708 60 720 63
rect 516 39 519 45
rect 525 39 528 45
rect 516 33 528 39
rect 516 27 519 33
rect 525 27 528 33
rect 516 21 528 27
rect 516 15 519 21
rect 525 15 528 21
rect 516 12 528 15
rect 612 45 624 48
rect 612 39 615 45
rect 621 39 624 45
rect 612 33 624 39
rect 612 27 615 33
rect 621 27 624 33
rect 612 21 624 27
rect 612 15 615 21
rect 621 15 624 21
rect 612 12 624 15
rect 636 45 648 48
rect 636 39 639 45
rect 645 39 648 45
rect 636 33 648 39
rect 636 27 639 33
rect 645 27 648 33
rect 636 21 648 27
rect 636 15 639 21
rect 645 15 648 21
rect 636 12 648 15
rect 732 45 744 255
rect 828 285 840 423
rect 900 429 912 519
rect 1044 477 1056 543
rect 1068 573 1080 576
rect 1068 567 1071 573
rect 1077 567 1080 573
rect 1068 561 1080 567
rect 1068 555 1071 561
rect 1077 555 1080 561
rect 1068 549 1080 555
rect 1068 543 1071 549
rect 1077 543 1080 549
rect 1068 540 1080 543
rect 1092 573 1104 576
rect 1092 567 1095 573
rect 1101 567 1104 573
rect 1092 561 1104 567
rect 1092 555 1095 561
rect 1101 555 1104 561
rect 1092 549 1104 555
rect 1092 543 1095 549
rect 1101 543 1104 549
rect 1044 471 1047 477
rect 1053 471 1056 477
rect 1044 465 1056 471
rect 1044 459 1047 465
rect 1053 459 1056 465
rect 1044 453 1056 459
rect 1044 447 1047 453
rect 1053 447 1056 453
rect 1044 444 1056 447
rect 1068 477 1080 480
rect 1068 471 1071 477
rect 1077 471 1080 477
rect 1068 465 1080 471
rect 1068 459 1071 465
rect 1077 459 1080 465
rect 1068 453 1080 459
rect 1068 447 1071 453
rect 1077 447 1080 453
rect 900 423 903 429
rect 909 423 912 429
rect 900 312 912 423
rect 1068 381 1080 447
rect 1092 477 1104 543
rect 1116 573 1128 576
rect 1116 567 1119 573
rect 1125 567 1128 573
rect 1116 561 1128 567
rect 1116 555 1119 561
rect 1125 555 1128 561
rect 1116 549 1128 555
rect 1116 543 1119 549
rect 1125 543 1128 549
rect 1116 540 1128 543
rect 1140 573 1152 576
rect 1140 567 1143 573
rect 1149 567 1152 573
rect 1140 561 1152 567
rect 1140 555 1143 561
rect 1149 555 1152 561
rect 1140 549 1152 555
rect 1140 543 1143 549
rect 1149 543 1152 549
rect 1116 525 1128 528
rect 1116 519 1119 525
rect 1125 519 1128 525
rect 1116 516 1128 519
rect 1092 471 1095 477
rect 1101 471 1104 477
rect 1092 465 1104 471
rect 1092 459 1095 465
rect 1101 459 1104 465
rect 1092 453 1104 459
rect 1092 447 1095 453
rect 1101 447 1104 453
rect 1092 444 1104 447
rect 1116 477 1128 480
rect 1116 471 1119 477
rect 1125 471 1128 477
rect 1116 465 1128 471
rect 1116 459 1119 465
rect 1125 459 1128 465
rect 1116 453 1128 459
rect 1116 447 1119 453
rect 1125 447 1128 453
rect 1092 429 1104 432
rect 1092 423 1095 429
rect 1101 423 1104 429
rect 1092 420 1104 423
rect 1068 375 1071 381
rect 1077 375 1080 381
rect 864 309 912 312
rect 864 303 867 309
rect 873 303 912 309
rect 864 300 912 303
rect 924 309 936 312
rect 924 303 927 309
rect 933 303 936 309
rect 924 300 936 303
rect 972 309 984 312
rect 972 303 975 309
rect 981 303 984 309
rect 972 300 984 303
rect 1020 309 1032 312
rect 1020 303 1023 309
rect 1029 303 1032 309
rect 1020 300 1032 303
rect 828 279 831 285
rect 837 279 840 285
rect 828 273 840 279
rect 828 267 831 273
rect 837 267 840 273
rect 828 261 840 267
rect 828 255 831 261
rect 837 255 840 261
rect 828 252 840 255
rect 852 285 864 288
rect 852 279 855 285
rect 861 279 864 285
rect 852 273 864 279
rect 852 267 855 273
rect 861 267 864 273
rect 852 261 864 267
rect 852 255 855 261
rect 861 255 864 261
rect 852 252 864 255
rect 876 285 888 288
rect 876 279 879 285
rect 885 279 888 285
rect 876 273 888 279
rect 876 267 879 273
rect 885 267 888 273
rect 876 261 888 267
rect 876 255 879 261
rect 885 255 888 261
rect 876 252 888 255
rect 900 285 912 300
rect 900 279 903 285
rect 909 279 912 285
rect 900 273 912 279
rect 900 267 903 273
rect 909 267 912 273
rect 900 261 912 267
rect 900 255 903 261
rect 909 255 912 261
rect 900 252 912 255
rect 1044 285 1056 288
rect 1044 279 1047 285
rect 1053 279 1056 285
rect 1044 273 1056 279
rect 1044 267 1047 273
rect 1053 267 1056 273
rect 1044 261 1056 267
rect 1044 255 1047 261
rect 1053 255 1056 261
rect 756 69 768 72
rect 756 63 759 69
rect 765 63 768 69
rect 756 60 768 63
rect 804 69 816 72
rect 804 63 807 69
rect 813 63 816 69
rect 804 60 816 63
rect 876 69 888 72
rect 876 63 879 69
rect 885 63 888 69
rect 876 60 888 63
rect 924 69 936 72
rect 924 63 927 69
rect 933 63 936 69
rect 924 60 936 63
rect 972 69 984 72
rect 972 63 975 69
rect 981 63 984 69
rect 972 60 984 63
rect 1020 69 1032 72
rect 1020 63 1023 69
rect 1029 63 1032 69
rect 1020 60 1032 63
rect 732 39 735 45
rect 741 39 744 45
rect 732 33 744 39
rect 732 27 735 33
rect 741 27 744 33
rect 732 21 744 27
rect 732 15 735 21
rect 741 15 744 21
rect 732 12 744 15
rect 828 45 840 48
rect 828 39 831 45
rect 837 39 840 45
rect 828 33 840 39
rect 828 27 831 33
rect 837 27 840 33
rect 828 21 840 27
rect 828 15 831 21
rect 837 15 840 21
rect 828 12 840 15
rect 852 45 864 48
rect 852 39 855 45
rect 861 39 864 45
rect 852 33 864 39
rect 852 27 855 33
rect 861 27 864 33
rect 852 21 864 27
rect 852 15 855 21
rect 861 15 864 21
rect 852 12 864 15
rect 1044 45 1056 255
rect 1068 285 1080 375
rect 1116 381 1128 447
rect 1140 477 1152 543
rect 1164 573 1176 576
rect 1164 567 1167 573
rect 1173 567 1176 573
rect 1164 561 1176 567
rect 1164 555 1167 561
rect 1173 555 1176 561
rect 1164 549 1176 555
rect 1164 543 1167 549
rect 1173 543 1176 549
rect 1164 540 1176 543
rect 1188 573 1200 576
rect 1188 567 1191 573
rect 1197 567 1200 573
rect 1188 561 1200 567
rect 1188 555 1191 561
rect 1197 555 1200 561
rect 1188 549 1200 555
rect 1188 543 1191 549
rect 1197 543 1200 549
rect 1164 525 1176 528
rect 1164 519 1167 525
rect 1173 519 1176 525
rect 1164 516 1176 519
rect 1140 471 1143 477
rect 1149 471 1152 477
rect 1140 465 1152 471
rect 1140 459 1143 465
rect 1149 459 1152 465
rect 1140 453 1152 459
rect 1140 447 1143 453
rect 1149 447 1152 453
rect 1140 444 1152 447
rect 1164 477 1176 504
rect 1164 471 1167 477
rect 1173 471 1176 477
rect 1164 465 1176 471
rect 1164 459 1167 465
rect 1173 459 1176 465
rect 1164 453 1176 459
rect 1164 447 1167 453
rect 1173 447 1176 453
rect 1140 429 1152 432
rect 1140 423 1143 429
rect 1149 423 1152 429
rect 1140 420 1152 423
rect 1116 375 1119 381
rect 1125 375 1128 381
rect 1092 309 1104 312
rect 1092 303 1095 309
rect 1101 303 1104 309
rect 1092 300 1104 303
rect 1068 279 1071 285
rect 1077 279 1080 285
rect 1068 273 1080 279
rect 1116 285 1128 375
rect 1164 381 1176 447
rect 1188 477 1200 543
rect 1212 573 1224 576
rect 1212 567 1215 573
rect 1221 567 1224 573
rect 1212 561 1224 567
rect 1212 555 1215 561
rect 1221 555 1224 561
rect 1212 549 1224 555
rect 1212 543 1215 549
rect 1221 543 1224 549
rect 1212 540 1224 543
rect 1236 573 1248 576
rect 1236 567 1239 573
rect 1245 567 1248 573
rect 1236 561 1248 567
rect 1236 555 1239 561
rect 1245 555 1248 561
rect 1236 549 1248 555
rect 1236 543 1239 549
rect 1245 543 1248 549
rect 1212 525 1224 528
rect 1212 519 1215 525
rect 1221 519 1224 525
rect 1212 516 1224 519
rect 1188 471 1191 477
rect 1197 471 1200 477
rect 1188 465 1200 471
rect 1188 459 1191 465
rect 1197 459 1200 465
rect 1188 453 1200 459
rect 1188 447 1191 453
rect 1197 447 1200 453
rect 1188 444 1200 447
rect 1212 477 1224 480
rect 1212 471 1215 477
rect 1221 471 1224 477
rect 1212 465 1224 471
rect 1212 459 1215 465
rect 1221 459 1224 465
rect 1212 453 1224 459
rect 1212 447 1215 453
rect 1221 447 1224 453
rect 1188 429 1200 432
rect 1188 423 1191 429
rect 1197 423 1200 429
rect 1188 420 1200 423
rect 1164 375 1167 381
rect 1173 375 1176 381
rect 1140 309 1152 312
rect 1140 303 1143 309
rect 1149 303 1152 309
rect 1140 300 1152 303
rect 1116 279 1119 285
rect 1125 279 1128 285
rect 1116 276 1128 279
rect 1164 285 1176 375
rect 1212 381 1224 447
rect 1236 477 1248 543
rect 1260 573 1272 576
rect 1260 567 1263 573
rect 1269 567 1272 573
rect 1260 561 1272 567
rect 1260 555 1263 561
rect 1269 555 1272 561
rect 1260 549 1272 555
rect 1260 543 1263 549
rect 1269 543 1272 549
rect 1260 540 1272 543
rect 1284 573 1296 576
rect 1284 567 1287 573
rect 1293 567 1296 573
rect 1284 561 1296 567
rect 1284 555 1287 561
rect 1293 555 1296 561
rect 1284 549 1296 555
rect 1284 543 1287 549
rect 1293 543 1296 549
rect 1284 540 1296 543
rect 1308 573 1320 576
rect 1308 567 1311 573
rect 1317 567 1320 573
rect 1308 561 1320 567
rect 1308 555 1311 561
rect 1317 555 1320 561
rect 1308 549 1320 555
rect 1308 543 1311 549
rect 1317 543 1320 549
rect 1236 471 1239 477
rect 1245 471 1248 477
rect 1236 465 1248 471
rect 1236 459 1239 465
rect 1245 459 1248 465
rect 1236 453 1248 459
rect 1236 447 1239 453
rect 1245 447 1248 453
rect 1236 444 1248 447
rect 1260 477 1272 480
rect 1260 471 1263 477
rect 1269 471 1272 477
rect 1260 465 1272 471
rect 1260 459 1263 465
rect 1269 459 1272 465
rect 1260 453 1272 459
rect 1260 447 1263 453
rect 1269 447 1272 453
rect 1236 429 1248 432
rect 1236 423 1239 429
rect 1245 423 1248 429
rect 1236 420 1248 423
rect 1212 375 1215 381
rect 1221 375 1224 381
rect 1188 309 1200 312
rect 1188 303 1191 309
rect 1197 303 1200 309
rect 1188 300 1200 303
rect 1164 279 1167 285
rect 1173 279 1176 285
rect 1164 276 1176 279
rect 1212 285 1224 375
rect 1260 381 1272 447
rect 1260 375 1263 381
rect 1269 375 1272 381
rect 1236 309 1248 312
rect 1236 303 1239 309
rect 1245 303 1248 309
rect 1236 300 1248 303
rect 1212 279 1215 285
rect 1221 279 1224 285
rect 1212 276 1224 279
rect 1260 285 1272 375
rect 1260 279 1263 285
rect 1269 279 1272 285
rect 1068 267 1071 273
rect 1077 267 1080 273
rect 1068 261 1080 267
rect 1260 273 1272 279
rect 1260 267 1263 273
rect 1269 267 1272 273
rect 1068 255 1071 261
rect 1077 255 1080 261
rect 1068 252 1080 255
rect 1092 261 1248 264
rect 1092 255 1095 261
rect 1101 255 1143 261
rect 1149 255 1191 261
rect 1197 255 1239 261
rect 1245 255 1248 261
rect 1092 252 1248 255
rect 1260 261 1272 267
rect 1260 255 1263 261
rect 1269 255 1272 261
rect 1260 252 1272 255
rect 1284 477 1296 480
rect 1284 471 1287 477
rect 1293 471 1296 477
rect 1284 465 1296 471
rect 1284 459 1287 465
rect 1293 459 1296 465
rect 1284 453 1296 459
rect 1284 447 1287 453
rect 1293 447 1296 453
rect 1284 288 1296 447
rect 1308 477 1320 543
rect 1332 573 1344 576
rect 1332 567 1335 573
rect 1341 567 1344 573
rect 1332 561 1344 567
rect 1332 555 1335 561
rect 1341 555 1344 561
rect 1332 549 1344 555
rect 1332 543 1335 549
rect 1341 543 1344 549
rect 1332 540 1344 543
rect 1356 573 1368 576
rect 1356 567 1359 573
rect 1365 567 1368 573
rect 1356 561 1368 567
rect 1356 555 1359 561
rect 1365 555 1368 561
rect 1356 549 1368 555
rect 1356 543 1359 549
rect 1365 543 1368 549
rect 1332 525 1344 528
rect 1332 519 1335 525
rect 1341 519 1344 525
rect 1332 516 1344 519
rect 1308 471 1311 477
rect 1317 471 1320 477
rect 1308 465 1320 471
rect 1308 459 1311 465
rect 1317 459 1320 465
rect 1308 453 1320 459
rect 1308 447 1311 453
rect 1317 447 1320 453
rect 1308 444 1320 447
rect 1332 477 1344 480
rect 1332 471 1335 477
rect 1341 471 1344 477
rect 1332 465 1344 471
rect 1332 459 1335 465
rect 1341 459 1344 465
rect 1332 453 1344 459
rect 1332 447 1335 453
rect 1341 447 1344 453
rect 1308 429 1320 432
rect 1308 423 1311 429
rect 1317 423 1320 429
rect 1308 420 1320 423
rect 1308 309 1320 312
rect 1308 303 1311 309
rect 1317 303 1320 309
rect 1308 300 1320 303
rect 1332 288 1344 447
rect 1356 477 1368 543
rect 1380 573 1392 576
rect 1380 567 1383 573
rect 1389 567 1392 573
rect 1380 561 1392 567
rect 1380 555 1383 561
rect 1389 555 1392 561
rect 1380 549 1392 555
rect 1380 543 1383 549
rect 1389 543 1392 549
rect 1380 540 1392 543
rect 1404 573 1416 576
rect 1404 567 1407 573
rect 1413 567 1416 573
rect 1404 561 1416 567
rect 1404 555 1407 561
rect 1413 555 1416 561
rect 1404 549 1416 555
rect 1404 543 1407 549
rect 1413 543 1416 549
rect 1356 471 1359 477
rect 1365 471 1368 477
rect 1356 465 1368 471
rect 1356 459 1359 465
rect 1365 459 1368 465
rect 1356 453 1368 459
rect 1356 447 1359 453
rect 1365 447 1368 453
rect 1356 444 1368 447
rect 1380 525 1392 528
rect 1380 519 1383 525
rect 1389 519 1392 525
rect 1380 477 1392 519
rect 1380 471 1383 477
rect 1389 471 1392 477
rect 1380 465 1392 471
rect 1380 459 1383 465
rect 1389 459 1392 465
rect 1380 453 1392 459
rect 1380 447 1383 453
rect 1389 447 1392 453
rect 1356 429 1368 432
rect 1356 423 1359 429
rect 1365 423 1368 429
rect 1356 420 1368 423
rect 1356 309 1368 312
rect 1356 303 1359 309
rect 1365 303 1368 309
rect 1356 300 1368 303
rect 1380 288 1392 447
rect 1404 477 1416 543
rect 1428 573 1440 576
rect 1428 567 1431 573
rect 1437 567 1440 573
rect 1428 561 1440 567
rect 1428 555 1431 561
rect 1437 555 1440 561
rect 1428 549 1440 555
rect 1428 543 1431 549
rect 1437 543 1440 549
rect 1428 540 1440 543
rect 1452 573 1464 576
rect 1452 567 1455 573
rect 1461 567 1464 573
rect 1452 561 1464 567
rect 1452 555 1455 561
rect 1461 555 1464 561
rect 1452 549 1464 555
rect 1452 543 1455 549
rect 1461 543 1464 549
rect 1428 525 1440 528
rect 1428 519 1431 525
rect 1437 519 1440 525
rect 1428 516 1440 519
rect 1404 471 1407 477
rect 1413 471 1416 477
rect 1404 465 1416 471
rect 1404 459 1407 465
rect 1413 459 1416 465
rect 1404 453 1416 459
rect 1404 447 1407 453
rect 1413 447 1416 453
rect 1404 444 1416 447
rect 1428 477 1440 480
rect 1428 471 1431 477
rect 1437 471 1440 477
rect 1428 465 1440 471
rect 1428 459 1431 465
rect 1437 459 1440 465
rect 1428 453 1440 459
rect 1428 447 1431 453
rect 1437 447 1440 453
rect 1404 429 1416 432
rect 1404 423 1407 429
rect 1413 423 1416 429
rect 1404 420 1416 423
rect 1404 309 1416 312
rect 1404 303 1407 309
rect 1413 303 1416 309
rect 1404 300 1416 303
rect 1428 288 1440 447
rect 1452 477 1464 543
rect 1476 573 1488 576
rect 1476 567 1479 573
rect 1485 567 1488 573
rect 1476 561 1488 567
rect 1476 555 1479 561
rect 1485 555 1488 561
rect 1476 549 1488 555
rect 1476 543 1479 549
rect 1485 543 1488 549
rect 1476 540 1488 543
rect 1452 471 1455 477
rect 1461 471 1464 477
rect 1452 465 1464 471
rect 1452 459 1455 465
rect 1461 459 1464 465
rect 1452 453 1464 459
rect 1452 447 1455 453
rect 1461 447 1464 453
rect 1452 444 1464 447
rect 1476 477 1488 480
rect 1476 471 1479 477
rect 1485 471 1488 477
rect 1476 465 1488 471
rect 1476 459 1479 465
rect 1485 459 1488 465
rect 1476 453 1488 459
rect 1476 447 1479 453
rect 1485 447 1488 453
rect 1452 429 1464 432
rect 1452 423 1455 429
rect 1461 423 1464 429
rect 1452 420 1464 423
rect 1452 309 1464 312
rect 1452 303 1455 309
rect 1461 303 1464 309
rect 1452 300 1464 303
rect 1476 288 1488 447
rect 1284 285 1488 288
rect 1284 279 1287 285
rect 1293 279 1335 285
rect 1341 279 1383 285
rect 1389 279 1431 285
rect 1437 279 1479 285
rect 1485 279 1488 285
rect 1284 276 1488 279
rect 1284 273 1296 276
rect 1284 267 1287 273
rect 1293 267 1296 273
rect 1284 261 1296 267
rect 1476 273 1488 276
rect 1476 267 1479 273
rect 1485 267 1488 273
rect 1284 255 1287 261
rect 1293 255 1296 261
rect 1284 252 1296 255
rect 1308 261 1464 264
rect 1308 255 1311 261
rect 1317 255 1359 261
rect 1365 255 1407 261
rect 1413 255 1455 261
rect 1461 255 1464 261
rect 1308 252 1464 255
rect 1476 261 1488 267
rect 1476 255 1479 261
rect 1485 255 1488 261
rect 1476 252 1488 255
rect 1092 69 1104 72
rect 1092 63 1095 69
rect 1101 63 1104 69
rect 1092 60 1104 63
rect 1116 48 1128 252
rect 1140 69 1152 72
rect 1140 63 1143 69
rect 1149 63 1152 69
rect 1140 60 1152 63
rect 1188 69 1200 72
rect 1188 63 1191 69
rect 1197 63 1200 69
rect 1188 60 1200 63
rect 1212 48 1224 252
rect 1308 237 1320 252
rect 1308 231 1311 237
rect 1317 231 1320 237
rect 1308 228 1320 231
rect 1356 237 1368 252
rect 1356 231 1359 237
rect 1365 231 1368 237
rect 1356 228 1368 231
rect 1404 237 1416 252
rect 1404 231 1407 237
rect 1413 231 1416 237
rect 1404 228 1416 231
rect 1452 237 1464 252
rect 1452 231 1455 237
rect 1461 231 1464 237
rect 1452 228 1464 231
rect 1524 213 1536 216
rect 1524 207 1527 213
rect 1533 207 1536 213
rect 1524 204 1536 207
rect 1236 69 1248 72
rect 1236 63 1239 69
rect 1245 63 1248 69
rect 1236 60 1248 63
rect 1044 39 1047 45
rect 1053 39 1056 45
rect 1044 33 1056 39
rect 1044 27 1047 33
rect 1053 27 1056 33
rect 1044 21 1056 27
rect 1044 15 1047 21
rect 1053 15 1056 21
rect 1044 12 1056 15
rect 1068 45 1080 48
rect 1068 39 1071 45
rect 1077 39 1080 45
rect 1068 33 1080 39
rect 1092 45 1152 48
rect 1092 39 1095 45
rect 1101 39 1143 45
rect 1149 39 1152 45
rect 1092 36 1152 39
rect 1164 45 1176 48
rect 1164 39 1167 45
rect 1173 39 1176 45
rect 1068 27 1071 33
rect 1077 27 1080 33
rect 1068 24 1080 27
rect 1164 33 1176 39
rect 1188 45 1248 48
rect 1188 39 1191 45
rect 1197 39 1239 45
rect 1245 39 1248 45
rect 1188 36 1248 39
rect 1260 45 1272 48
rect 1260 39 1263 45
rect 1269 39 1272 45
rect 1164 27 1167 33
rect 1173 27 1176 33
rect 1164 24 1176 27
rect 1260 33 1272 39
rect 1260 27 1263 33
rect 1269 27 1272 33
rect 1260 24 1272 27
rect 1068 21 1272 24
rect 1068 15 1071 21
rect 1077 15 1119 21
rect 1125 15 1167 21
rect 1173 15 1215 21
rect 1221 15 1263 21
rect 1269 15 1272 21
rect 1068 12 1272 15
<< via2 >>
rect -9 567 -3 573
rect -9 555 -3 561
rect -9 543 -3 549
rect -9 495 -3 501
rect -9 447 -3 453
rect -33 399 -27 405
rect -33 351 -27 357
rect 39 567 45 573
rect 39 555 45 561
rect 39 543 45 549
rect 39 519 45 525
rect 15 471 21 477
rect 39 447 45 453
rect 15 423 21 429
rect 87 567 93 573
rect 87 555 93 561
rect 87 543 93 549
rect 87 519 93 525
rect 63 471 69 477
rect 87 447 93 453
rect 63 423 69 429
rect 135 567 141 573
rect 135 555 141 561
rect 135 543 141 549
rect 135 519 141 525
rect 111 471 117 477
rect 135 447 141 453
rect 111 423 117 429
rect 183 567 189 573
rect 183 555 189 561
rect 183 543 189 549
rect 207 567 213 573
rect 207 555 213 561
rect 207 543 213 549
rect 231 519 237 525
rect 159 471 165 477
rect 183 447 189 453
rect 159 423 165 429
rect 207 447 213 453
rect -57 207 -51 213
rect -9 183 -3 189
rect 39 183 45 189
rect 87 183 93 189
rect 39 159 45 165
rect 15 63 21 69
rect -9 39 -3 45
rect -9 27 -3 33
rect -9 15 -3 21
rect 63 63 69 69
rect 135 183 141 189
rect 303 567 309 573
rect 303 555 309 561
rect 303 543 309 549
rect 279 519 285 525
rect 327 519 333 525
rect 255 471 261 477
rect 303 447 309 453
rect 399 567 405 573
rect 399 555 405 561
rect 399 543 405 549
rect 423 567 429 573
rect 423 555 429 561
rect 423 543 429 549
rect 375 519 381 525
rect 351 471 357 477
rect 399 447 405 453
rect 231 423 237 429
rect 279 423 285 429
rect 327 423 333 429
rect 375 423 381 429
rect 231 303 237 309
rect 279 303 285 309
rect 327 303 333 309
rect 375 303 381 309
rect 183 183 189 189
rect 135 159 141 165
rect 111 63 117 69
rect 255 159 261 165
rect 159 63 165 69
rect 231 63 237 69
rect 183 39 189 45
rect 183 27 189 33
rect 183 15 189 21
rect 207 39 213 45
rect 207 27 213 33
rect 207 15 213 21
rect 423 447 429 453
rect 519 567 525 573
rect 519 555 525 561
rect 519 543 525 549
rect 519 519 525 525
rect 471 471 477 477
rect 519 447 525 453
rect 615 567 621 573
rect 615 555 621 561
rect 615 543 621 549
rect 639 567 645 573
rect 639 555 645 561
rect 639 543 645 549
rect 567 471 573 477
rect 615 447 621 453
rect 447 423 453 429
rect 495 423 501 429
rect 543 423 549 429
rect 591 423 597 429
rect 423 303 429 309
rect 447 303 453 309
rect 495 303 501 309
rect 543 303 549 309
rect 591 303 597 309
rect 303 135 309 141
rect 279 63 285 69
rect 351 159 357 165
rect 327 63 333 69
rect 639 423 645 429
rect 663 423 669 429
rect 711 423 717 429
rect 759 423 765 429
rect 807 423 813 429
rect 663 303 669 309
rect 711 303 717 309
rect 759 303 765 309
rect 807 303 813 309
rect 519 111 525 117
rect 375 63 381 69
rect 447 63 453 69
rect 495 63 501 69
rect 399 39 405 45
rect 399 27 405 33
rect 399 15 405 21
rect 423 39 429 45
rect 423 27 429 33
rect 423 15 429 21
rect 543 63 549 69
rect 591 63 597 69
rect 663 63 669 69
rect 711 63 717 69
rect 615 39 621 45
rect 615 27 621 33
rect 615 15 621 21
rect 639 39 645 45
rect 639 27 645 33
rect 639 15 645 21
rect 1071 567 1077 573
rect 1071 555 1077 561
rect 1071 543 1077 549
rect 1119 567 1125 573
rect 1119 555 1125 561
rect 1119 543 1125 549
rect 1119 519 1125 525
rect 1095 471 1101 477
rect 1095 423 1101 429
rect 1071 375 1077 381
rect 927 303 933 309
rect 975 303 981 309
rect 1023 303 1029 309
rect 759 63 765 69
rect 807 63 813 69
rect 879 63 885 69
rect 927 63 933 69
rect 975 63 981 69
rect 1023 63 1029 69
rect 831 39 837 45
rect 831 27 837 33
rect 831 15 837 21
rect 855 39 861 45
rect 855 27 861 33
rect 855 15 861 21
rect 1167 567 1173 573
rect 1167 555 1173 561
rect 1167 543 1173 549
rect 1167 519 1173 525
rect 1143 471 1149 477
rect 1143 423 1149 429
rect 1119 375 1125 381
rect 1095 303 1101 309
rect 1071 279 1077 285
rect 1215 567 1221 573
rect 1215 555 1221 561
rect 1215 543 1221 549
rect 1215 519 1221 525
rect 1191 471 1197 477
rect 1191 423 1197 429
rect 1167 375 1173 381
rect 1143 303 1149 309
rect 1119 279 1125 285
rect 1263 567 1269 573
rect 1263 555 1269 561
rect 1263 543 1269 549
rect 1287 567 1293 573
rect 1287 555 1293 561
rect 1287 543 1293 549
rect 1239 471 1245 477
rect 1239 423 1245 429
rect 1215 375 1221 381
rect 1191 303 1197 309
rect 1167 279 1173 285
rect 1263 375 1269 381
rect 1239 303 1245 309
rect 1215 279 1221 285
rect 1263 279 1269 285
rect 1335 567 1341 573
rect 1335 555 1341 561
rect 1335 543 1341 549
rect 1335 519 1341 525
rect 1311 471 1317 477
rect 1311 423 1317 429
rect 1311 303 1317 309
rect 1383 567 1389 573
rect 1383 555 1389 561
rect 1383 543 1389 549
rect 1359 471 1365 477
rect 1383 519 1389 525
rect 1359 423 1365 429
rect 1359 303 1365 309
rect 1431 567 1437 573
rect 1431 555 1437 561
rect 1431 543 1437 549
rect 1431 519 1437 525
rect 1407 471 1413 477
rect 1407 423 1413 429
rect 1407 303 1413 309
rect 1479 567 1485 573
rect 1479 555 1485 561
rect 1479 543 1485 549
rect 1455 471 1461 477
rect 1455 423 1461 429
rect 1455 303 1461 309
rect 1095 63 1101 69
rect 1143 63 1149 69
rect 1191 63 1197 69
rect 1311 231 1317 237
rect 1359 231 1365 237
rect 1407 231 1413 237
rect 1455 231 1461 237
rect 1527 207 1533 213
rect 1239 63 1245 69
rect 1071 39 1077 45
rect 1167 39 1173 45
rect 1071 27 1077 33
rect 1263 39 1269 45
rect 1167 27 1173 33
rect 1263 27 1269 33
rect 1071 15 1077 21
rect 1167 15 1173 21
rect 1263 15 1269 21
<< metal3 >>
rect -60 573 1536 576
rect -60 567 -9 573
rect -3 567 39 573
rect 45 567 87 573
rect 93 567 135 573
rect 141 567 183 573
rect 189 567 207 573
rect 213 567 303 573
rect 309 567 399 573
rect 405 567 423 573
rect 429 567 519 573
rect 525 567 615 573
rect 621 567 639 573
rect 645 567 1071 573
rect 1077 567 1119 573
rect 1125 567 1167 573
rect 1173 567 1215 573
rect 1221 567 1263 573
rect 1269 567 1287 573
rect 1293 567 1335 573
rect 1341 567 1383 573
rect 1389 567 1431 573
rect 1437 567 1479 573
rect 1485 567 1536 573
rect -60 561 1536 567
rect -60 555 -9 561
rect -3 555 39 561
rect 45 555 87 561
rect 93 555 135 561
rect 141 555 183 561
rect 189 555 207 561
rect 213 555 303 561
rect 309 555 399 561
rect 405 555 423 561
rect 429 555 519 561
rect 525 555 615 561
rect 621 555 639 561
rect 645 555 1071 561
rect 1077 555 1119 561
rect 1125 555 1167 561
rect 1173 555 1215 561
rect 1221 555 1263 561
rect 1269 555 1287 561
rect 1293 555 1335 561
rect 1341 555 1383 561
rect 1389 555 1431 561
rect 1437 555 1479 561
rect 1485 555 1536 561
rect -60 549 1536 555
rect -60 543 -9 549
rect -3 543 39 549
rect 45 543 87 549
rect 93 543 135 549
rect 141 543 183 549
rect 189 543 207 549
rect 213 543 303 549
rect 309 543 399 549
rect 405 543 423 549
rect 429 543 519 549
rect 525 543 615 549
rect 621 543 639 549
rect 645 543 1071 549
rect 1077 543 1119 549
rect 1125 543 1167 549
rect 1173 543 1215 549
rect 1221 543 1263 549
rect 1269 543 1287 549
rect 1293 543 1335 549
rect 1341 543 1383 549
rect 1389 543 1431 549
rect 1437 543 1479 549
rect 1485 543 1536 549
rect -60 540 1536 543
rect -24 525 1056 528
rect -24 519 39 525
rect 45 519 87 525
rect 93 519 135 525
rect 141 519 231 525
rect 237 519 279 525
rect 285 519 303 525
rect 309 519 327 525
rect 333 519 375 525
rect 381 519 519 525
rect 525 519 855 525
rect 861 519 1056 525
rect -24 516 1056 519
rect 1068 525 1488 528
rect 1068 519 1119 525
rect 1125 519 1167 525
rect 1173 519 1215 525
rect 1221 519 1335 525
rect 1341 519 1383 525
rect 1389 519 1431 525
rect 1437 519 1488 525
rect 1068 516 1488 519
rect -60 501 1512 504
rect -60 495 -9 501
rect -3 495 1512 501
rect -60 492 1512 495
rect 12 477 168 480
rect 12 471 15 477
rect 21 471 63 477
rect 69 471 111 477
rect 117 471 159 477
rect 165 471 168 477
rect 12 468 168 471
rect 252 477 360 480
rect 252 471 255 477
rect 261 471 351 477
rect 357 471 360 477
rect 252 468 360 471
rect 468 477 576 480
rect 468 471 471 477
rect 477 471 567 477
rect 573 471 576 477
rect 468 468 576 471
rect 1092 477 1248 480
rect 1092 471 1095 477
rect 1101 471 1143 477
rect 1149 471 1191 477
rect 1197 471 1239 477
rect 1245 471 1248 477
rect 1092 468 1248 471
rect 1308 477 1464 480
rect 1308 471 1311 477
rect 1317 471 1359 477
rect 1365 471 1407 477
rect 1413 471 1455 477
rect 1461 471 1464 477
rect 1308 468 1464 471
rect -12 453 192 456
rect -12 447 -9 453
rect -3 447 39 453
rect 45 447 87 453
rect 93 447 135 453
rect 141 447 183 453
rect 189 447 192 453
rect -12 444 192 447
rect 204 453 408 456
rect 204 447 207 453
rect 213 447 303 453
rect 309 447 399 453
rect 405 447 408 453
rect 204 444 408 447
rect 420 453 624 456
rect 420 447 423 453
rect 429 447 519 453
rect 525 447 615 453
rect 621 447 624 453
rect 420 444 624 447
rect -24 429 1488 432
rect -24 423 15 429
rect 21 423 63 429
rect 69 423 111 429
rect 117 423 159 429
rect 165 423 231 429
rect 237 423 279 429
rect 285 423 327 429
rect 333 423 375 429
rect 381 423 447 429
rect 453 423 495 429
rect 501 423 543 429
rect 549 423 591 429
rect 597 423 639 429
rect 645 423 663 429
rect 669 423 711 429
rect 717 423 759 429
rect 765 423 807 429
rect 813 423 1095 429
rect 1101 423 1143 429
rect 1149 423 1191 429
rect 1197 423 1239 429
rect 1245 423 1311 429
rect 1317 423 1359 429
rect 1365 423 1407 429
rect 1413 423 1455 429
rect 1461 423 1488 429
rect -24 420 1488 423
rect -36 405 1512 408
rect -36 399 -33 405
rect -27 399 1512 405
rect -36 396 1512 399
rect -36 381 1536 384
rect -36 375 1071 381
rect 1077 375 1119 381
rect 1125 375 1167 381
rect 1173 375 1215 381
rect 1221 375 1263 381
rect 1269 375 1536 381
rect -36 372 1536 375
rect -48 357 1512 360
rect -48 351 -33 357
rect -27 351 1512 357
rect -48 348 1512 351
rect 216 309 1500 312
rect 216 303 231 309
rect 237 303 279 309
rect 285 303 327 309
rect 333 303 375 309
rect 381 303 423 309
rect 429 303 447 309
rect 453 303 495 309
rect 501 303 543 309
rect 549 303 591 309
rect 597 303 663 309
rect 669 303 711 309
rect 717 303 759 309
rect 765 303 807 309
rect 813 303 927 309
rect 933 303 975 309
rect 981 303 1023 309
rect 1029 303 1095 309
rect 1101 303 1143 309
rect 1149 303 1191 309
rect 1197 303 1239 309
rect 1245 303 1311 309
rect 1317 303 1359 309
rect 1365 303 1407 309
rect 1413 303 1455 309
rect 1461 303 1500 309
rect 216 300 1500 303
rect 852 285 864 288
rect 852 279 855 285
rect 861 279 864 285
rect 852 273 864 279
rect 852 267 855 273
rect 861 267 864 273
rect 852 261 864 267
rect 852 255 855 261
rect 861 255 864 261
rect 852 252 864 255
rect 876 285 888 288
rect 876 279 879 285
rect 885 279 888 285
rect 876 273 888 279
rect 1068 285 1272 288
rect 1068 279 1071 285
rect 1077 279 1119 285
rect 1125 279 1167 285
rect 1173 279 1215 285
rect 1221 279 1263 285
rect 1269 279 1272 285
rect 1068 276 1272 279
rect 876 267 879 273
rect 885 267 888 273
rect 876 261 888 267
rect 876 255 879 261
rect 885 255 888 261
rect 876 252 888 255
rect -24 237 1536 240
rect -24 231 1311 237
rect 1317 231 1359 237
rect 1365 231 1407 237
rect 1413 231 1455 237
rect 1461 231 1536 237
rect -24 228 1536 231
rect -60 213 1536 216
rect -60 207 -57 213
rect -51 207 1527 213
rect 1533 207 1536 213
rect -60 204 1536 207
rect -24 189 1500 192
rect -24 183 -9 189
rect -3 183 15 189
rect 21 183 39 189
rect 45 183 63 189
rect 69 183 87 189
rect 93 183 111 189
rect 117 183 135 189
rect 141 183 159 189
rect 165 183 183 189
rect 189 183 231 189
rect 237 183 375 189
rect 381 183 1500 189
rect -24 180 1500 183
rect -24 165 1500 168
rect -24 159 39 165
rect 45 159 135 165
rect 141 159 255 165
rect 261 159 351 165
rect 357 159 1500 165
rect -24 156 1500 159
rect -24 141 1500 144
rect -24 135 303 141
rect 309 135 1500 141
rect -24 132 1500 135
rect -24 117 1500 120
rect -24 111 279 117
rect 285 111 327 117
rect 333 111 447 117
rect 453 111 495 117
rect 501 111 519 117
rect 525 111 543 117
rect 549 111 591 117
rect 597 111 663 117
rect 669 111 711 117
rect 717 111 759 117
rect 765 111 807 117
rect 813 111 879 117
rect 885 111 927 117
rect 933 111 975 117
rect 981 111 1023 117
rect 1029 111 1095 117
rect 1101 111 1143 117
rect 1149 111 1191 117
rect 1197 111 1239 117
rect 1245 111 1500 117
rect -24 108 1500 111
rect 12 69 24 72
rect 12 63 15 69
rect 21 63 24 69
rect 12 60 24 63
rect 60 69 72 72
rect 60 63 63 69
rect 69 63 72 69
rect 60 60 72 63
rect 108 69 120 72
rect 108 63 111 69
rect 117 63 120 69
rect 108 60 120 63
rect 156 69 168 72
rect 156 63 159 69
rect 165 63 168 69
rect 156 60 168 63
rect 228 69 240 72
rect 228 63 231 69
rect 237 63 240 69
rect 228 60 240 63
rect 276 69 288 72
rect 276 63 279 69
rect 285 63 288 69
rect 276 60 288 63
rect 324 69 336 72
rect 324 63 327 69
rect 333 63 336 69
rect 324 60 336 63
rect 372 69 384 72
rect 372 63 375 69
rect 381 63 384 69
rect 372 60 384 63
rect 444 69 456 72
rect 444 63 447 69
rect 453 63 456 69
rect 444 60 456 63
rect 492 69 504 72
rect 492 63 495 69
rect 501 63 504 69
rect 492 60 504 63
rect 540 69 552 72
rect 540 63 543 69
rect 549 63 552 69
rect 540 60 552 63
rect 588 69 600 72
rect 588 63 591 69
rect 597 63 600 69
rect 588 60 600 63
rect 660 69 672 72
rect 660 63 663 69
rect 669 63 672 69
rect 660 60 672 63
rect 708 69 720 72
rect 708 63 711 69
rect 717 63 720 69
rect 708 60 720 63
rect 756 69 768 72
rect 756 63 759 69
rect 765 63 768 69
rect 756 60 768 63
rect 804 69 816 72
rect 804 63 807 69
rect 813 63 816 69
rect 804 60 816 63
rect 876 69 888 72
rect 876 63 879 69
rect 885 63 888 69
rect 876 60 888 63
rect 924 69 936 72
rect 924 63 927 69
rect 933 63 936 69
rect 924 60 936 63
rect 972 69 984 72
rect 972 63 975 69
rect 981 63 984 69
rect 972 60 984 63
rect 1020 69 1032 72
rect 1020 63 1023 69
rect 1029 63 1032 69
rect 1020 60 1032 63
rect 1092 69 1104 72
rect 1092 63 1095 69
rect 1101 63 1104 69
rect 1092 60 1104 63
rect 1140 69 1152 72
rect 1140 63 1143 69
rect 1149 63 1152 69
rect 1140 60 1152 63
rect 1188 69 1200 72
rect 1188 63 1191 69
rect 1197 63 1200 69
rect 1188 60 1200 63
rect 1236 69 1248 72
rect 1236 63 1239 69
rect 1245 63 1248 69
rect 1236 60 1248 63
rect -60 45 1536 48
rect -60 39 -9 45
rect -3 39 183 45
rect 189 39 207 45
rect 213 39 399 45
rect 405 39 423 45
rect 429 39 615 45
rect 621 39 639 45
rect 645 39 831 45
rect 837 39 855 45
rect 861 39 1071 45
rect 1077 39 1167 45
rect 1173 39 1263 45
rect 1269 39 1536 45
rect -60 33 1536 39
rect -60 27 -9 33
rect -3 27 183 33
rect 189 27 207 33
rect 213 27 399 33
rect 405 27 423 33
rect 429 27 615 33
rect 621 27 639 33
rect 645 27 831 33
rect 837 27 855 33
rect 861 27 1071 33
rect 1077 27 1167 33
rect 1173 27 1263 33
rect 1269 27 1536 33
rect -60 21 1536 27
rect -60 15 -9 21
rect -3 15 183 21
rect 189 15 207 21
rect 213 15 399 21
rect 405 15 423 21
rect 429 15 615 21
rect 621 15 639 21
rect 645 15 831 21
rect 837 15 855 21
rect 861 15 1071 21
rect 1077 15 1167 21
rect 1173 15 1263 21
rect 1269 15 1536 21
rect -60 12 1536 15
<< via3 >>
rect 303 519 309 525
rect 855 519 861 525
rect 303 447 309 453
rect 855 279 861 285
rect 855 267 861 273
rect 855 255 861 261
rect 879 279 885 285
rect 879 267 885 273
rect 879 255 885 261
rect 15 183 21 189
rect 63 183 69 189
rect 111 183 117 189
rect 159 183 165 189
rect 231 183 237 189
rect 375 183 381 189
rect 279 111 285 117
rect 327 111 333 117
rect 447 111 453 117
rect 495 111 501 117
rect 543 111 549 117
rect 591 111 597 117
rect 663 111 669 117
rect 711 111 717 117
rect 759 111 765 117
rect 807 111 813 117
rect 879 111 885 117
rect 927 111 933 117
rect 975 111 981 117
rect 1023 111 1029 117
rect 1095 111 1101 117
rect 1143 111 1149 117
rect 1191 111 1197 117
rect 1239 111 1245 117
rect 15 63 21 69
rect 63 63 69 69
rect 111 63 117 69
rect 159 63 165 69
rect 231 63 237 69
rect 279 63 285 69
rect 327 63 333 69
rect 375 63 381 69
rect 447 63 453 69
rect 495 63 501 69
rect 543 63 549 69
rect 591 63 597 69
rect 663 63 669 69
rect 711 63 717 69
rect 759 63 765 69
rect 807 63 813 69
rect 879 63 885 69
rect 927 63 933 69
rect 975 63 981 69
rect 1023 63 1029 69
rect 1095 63 1101 69
rect 1143 63 1149 69
rect 1191 63 1197 69
rect 1239 63 1245 69
<< metal4 >>
rect 852 552 864 576
rect 300 525 312 528
rect 300 519 303 525
rect 309 519 312 525
rect 300 453 312 519
rect 300 447 303 453
rect 309 447 312 453
rect 300 444 312 447
rect 852 525 864 528
rect 852 519 855 525
rect 861 519 864 525
rect 192 396 204 408
rect 408 396 420 408
rect 624 396 636 408
rect 192 324 204 360
rect 408 324 420 360
rect 624 324 636 360
rect 852 285 864 519
rect 852 279 855 285
rect 861 279 864 285
rect 852 273 864 279
rect 852 267 855 273
rect 861 267 864 273
rect 852 261 864 267
rect 852 255 855 261
rect 861 255 864 261
rect 852 252 864 255
rect 876 285 888 288
rect 876 279 879 285
rect 885 279 888 285
rect 876 273 888 279
rect 876 267 879 273
rect 885 267 888 273
rect 876 261 888 267
rect 876 255 879 261
rect 885 255 888 261
rect 12 204 24 216
rect 60 204 72 216
rect 108 204 120 216
rect 156 204 168 216
rect 228 204 240 216
rect 276 204 288 216
rect 324 204 336 216
rect 372 204 384 216
rect 444 204 456 216
rect 492 204 504 216
rect 540 204 552 216
rect 588 204 600 216
rect 660 204 672 216
rect 708 204 720 216
rect 756 204 768 216
rect 804 204 816 216
rect 12 189 24 192
rect 12 183 15 189
rect 21 183 24 189
rect 12 69 24 183
rect 12 63 15 69
rect 21 63 24 69
rect 12 60 24 63
rect 60 189 72 192
rect 60 183 63 189
rect 69 183 72 189
rect 60 69 72 183
rect 60 63 63 69
rect 69 63 72 69
rect 60 60 72 63
rect 108 189 120 192
rect 108 183 111 189
rect 117 183 120 189
rect 108 69 120 183
rect 108 63 111 69
rect 117 63 120 69
rect 108 60 120 63
rect 156 189 168 192
rect 156 183 159 189
rect 165 183 168 189
rect 156 69 168 183
rect 156 63 159 69
rect 165 63 168 69
rect 156 60 168 63
rect 228 189 240 192
rect 228 183 231 189
rect 237 183 240 189
rect 228 69 240 183
rect 372 189 384 192
rect 372 183 375 189
rect 381 183 384 189
rect 228 63 231 69
rect 237 63 240 69
rect 228 60 240 63
rect 276 117 288 120
rect 276 111 279 117
rect 285 111 288 117
rect 276 69 288 111
rect 276 63 279 69
rect 285 63 288 69
rect 276 60 288 63
rect 324 117 336 120
rect 324 111 327 117
rect 333 111 336 117
rect 324 69 336 111
rect 324 63 327 69
rect 333 63 336 69
rect 324 60 336 63
rect 372 69 384 183
rect 372 63 375 69
rect 381 63 384 69
rect 372 60 384 63
rect 444 117 456 120
rect 444 111 447 117
rect 453 111 456 117
rect 444 69 456 111
rect 444 63 447 69
rect 453 63 456 69
rect 444 60 456 63
rect 492 117 504 120
rect 492 111 495 117
rect 501 111 504 117
rect 492 69 504 111
rect 492 63 495 69
rect 501 63 504 69
rect 492 60 504 63
rect 540 117 552 120
rect 540 111 543 117
rect 549 111 552 117
rect 540 69 552 111
rect 540 63 543 69
rect 549 63 552 69
rect 540 60 552 63
rect 588 117 600 120
rect 588 111 591 117
rect 597 111 600 117
rect 588 69 600 111
rect 588 63 591 69
rect 597 63 600 69
rect 588 60 600 63
rect 660 117 672 120
rect 660 111 663 117
rect 669 111 672 117
rect 660 69 672 111
rect 660 63 663 69
rect 669 63 672 69
rect 660 60 672 63
rect 708 117 720 120
rect 708 111 711 117
rect 717 111 720 117
rect 708 69 720 111
rect 708 63 711 69
rect 717 63 720 69
rect 708 60 720 63
rect 756 117 768 120
rect 756 111 759 117
rect 765 111 768 117
rect 756 69 768 111
rect 756 63 759 69
rect 765 63 768 69
rect 756 60 768 63
rect 804 117 816 120
rect 804 111 807 117
rect 813 111 816 117
rect 804 69 816 111
rect 804 63 807 69
rect 813 63 816 69
rect 804 60 816 63
rect 876 117 888 255
rect 924 204 936 216
rect 972 204 984 216
rect 1020 204 1032 216
rect 1092 204 1104 216
rect 1140 204 1152 216
rect 1188 204 1200 216
rect 1236 204 1248 216
rect 876 111 879 117
rect 885 111 888 117
rect 876 69 888 111
rect 876 63 879 69
rect 885 63 888 69
rect 876 60 888 63
rect 924 117 936 120
rect 924 111 927 117
rect 933 111 936 117
rect 924 69 936 111
rect 924 63 927 69
rect 933 63 936 69
rect 924 60 936 63
rect 972 117 984 120
rect 972 111 975 117
rect 981 111 984 117
rect 972 69 984 111
rect 972 63 975 69
rect 981 63 984 69
rect 972 60 984 63
rect 1020 117 1032 120
rect 1020 111 1023 117
rect 1029 111 1032 117
rect 1020 69 1032 111
rect 1020 63 1023 69
rect 1029 63 1032 69
rect 1020 60 1032 63
rect 1092 117 1104 120
rect 1092 111 1095 117
rect 1101 111 1104 117
rect 1092 69 1104 111
rect 1092 63 1095 69
rect 1101 63 1104 69
rect 1092 60 1104 63
rect 1140 117 1152 120
rect 1140 111 1143 117
rect 1149 111 1152 117
rect 1140 69 1152 111
rect 1140 63 1143 69
rect 1149 63 1152 69
rect 1140 60 1152 63
rect 1188 117 1200 120
rect 1188 111 1191 117
rect 1197 111 1200 117
rect 1188 69 1200 111
rect 1188 63 1191 69
rect 1197 63 1200 69
rect 1188 60 1200 63
rect 1236 117 1248 120
rect 1236 111 1239 117
rect 1245 111 1248 117
rect 1236 69 1248 111
rect 1236 63 1239 69
rect 1245 63 1248 69
rect 1236 60 1248 63
<< labels >>
rlabel metal3 1524 228 1536 240 0 iq
port 1 nsew
rlabel metal3 1524 372 1536 384 0 gp
port 2 nsew
rlabel metal3 -24 108 -12 120 0 bn
rlabel metal3 -24 132 -12 144 0 bn0
rlabel metal3 -24 156 -12 168 0 y
rlabel metal3 -24 180 -12 192 0 x
rlabel metal2 900 312 912 324 0 s
rlabel metal3 -60 540 -48 576 0 vdd
port 3 nsew
rlabel metal3 -60 12 -48 48 0 vss
port 4 nsew
rlabel metal3 -24 516 -12 528 0 bpa
rlabel metal3 -24 420 -12 432 0 bpb
rlabel metal3 1524 540 1536 576 0 vdd
port 3 nsew
<< end >>
