magic
tech gf180mcuC
timestamp 1697197950
<< nwell >>
rect -42 -30 102 102
rect 126 -30 270 102
rect -42 -186 102 -54
rect 126 -186 270 -54
rect -42 -342 102 -210
<< nmos >>
rect 168 -300 228 -264
<< mvpmos >>
rect 0 12 60 48
rect 168 12 228 48
rect 0 -132 60 -96
rect 168 -132 228 -96
rect 0 -300 60 -264
<< ndiff >>
rect 156 -267 168 -264
rect 156 -273 159 -267
rect 165 -273 168 -267
rect 156 -279 168 -273
rect 156 -285 159 -279
rect 165 -285 168 -279
rect 156 -291 168 -285
rect 156 -297 159 -291
rect 165 -297 168 -291
rect 156 -300 168 -297
rect 228 -267 240 -264
rect 228 -273 231 -267
rect 237 -273 240 -267
rect 228 -279 240 -273
rect 228 -285 231 -279
rect 237 -285 240 -279
rect 228 -291 240 -285
rect 228 -297 231 -291
rect 237 -297 240 -291
rect 228 -300 240 -297
<< mvpdiff >>
rect -12 45 0 48
rect -12 39 -9 45
rect -3 39 0 45
rect -12 33 0 39
rect -12 27 -9 33
rect -3 27 0 33
rect -12 21 0 27
rect -12 15 -9 21
rect -3 15 0 21
rect -12 12 0 15
rect 60 45 72 48
rect 60 39 63 45
rect 69 39 72 45
rect 60 33 72 39
rect 60 27 63 33
rect 69 27 72 33
rect 60 21 72 27
rect 60 15 63 21
rect 69 15 72 21
rect 60 12 72 15
rect 156 45 168 48
rect 156 39 159 45
rect 165 39 168 45
rect 156 33 168 39
rect 156 27 159 33
rect 165 27 168 33
rect 156 21 168 27
rect 156 15 159 21
rect 165 15 168 21
rect 156 12 168 15
rect 228 45 240 48
rect 228 39 231 45
rect 237 39 240 45
rect 228 33 240 39
rect 228 27 231 33
rect 237 27 240 33
rect 228 21 240 27
rect 228 15 231 21
rect 237 15 240 21
rect 228 12 240 15
rect -12 -99 0 -96
rect -12 -105 -9 -99
rect -3 -105 0 -99
rect -12 -111 0 -105
rect -12 -117 -9 -111
rect -3 -117 0 -111
rect -12 -123 0 -117
rect -12 -129 -9 -123
rect -3 -129 0 -123
rect -12 -132 0 -129
rect 60 -99 72 -96
rect 60 -105 63 -99
rect 69 -105 72 -99
rect 60 -111 72 -105
rect 60 -117 63 -111
rect 69 -117 72 -111
rect 60 -123 72 -117
rect 60 -129 63 -123
rect 69 -129 72 -123
rect 60 -132 72 -129
rect 156 -99 168 -96
rect 156 -105 159 -99
rect 165 -105 168 -99
rect 156 -111 168 -105
rect 156 -117 159 -111
rect 165 -117 168 -111
rect 156 -123 168 -117
rect 156 -129 159 -123
rect 165 -129 168 -123
rect 156 -132 168 -129
rect 228 -99 240 -96
rect 228 -105 231 -99
rect 237 -105 240 -99
rect 228 -111 240 -105
rect 228 -117 231 -111
rect 237 -117 240 -111
rect 228 -123 240 -117
rect 228 -129 231 -123
rect 237 -129 240 -123
rect 228 -132 240 -129
rect -12 -267 0 -264
rect -12 -273 -9 -267
rect -3 -273 0 -267
rect -12 -279 0 -273
rect -12 -285 -9 -279
rect -3 -285 0 -279
rect -12 -291 0 -285
rect -12 -297 -9 -291
rect -3 -297 0 -291
rect -12 -300 0 -297
rect 60 -267 72 -264
rect 60 -273 63 -267
rect 69 -273 72 -267
rect 60 -279 72 -273
rect 60 -285 63 -279
rect 69 -285 72 -279
rect 60 -291 72 -285
rect 60 -297 63 -291
rect 69 -297 72 -291
rect 60 -300 72 -297
<< ndiffc >>
rect 159 -273 165 -267
rect 159 -285 165 -279
rect 159 -297 165 -291
rect 231 -273 237 -267
rect 231 -285 237 -279
rect 231 -297 237 -291
<< mvpdiffc >>
rect -9 39 -3 45
rect -9 27 -3 33
rect -9 15 -3 21
rect 63 39 69 45
rect 63 27 69 33
rect 63 15 69 21
rect 159 39 165 45
rect 159 27 165 33
rect 159 15 165 21
rect 231 39 237 45
rect 231 27 237 33
rect 231 15 237 21
rect -9 -105 -3 -99
rect -9 -117 -3 -111
rect -9 -129 -3 -123
rect 63 -105 69 -99
rect 63 -117 69 -111
rect 63 -129 69 -123
rect 159 -105 165 -99
rect 159 -117 165 -111
rect 159 -129 165 -123
rect 231 -105 237 -99
rect 231 -117 237 -111
rect 231 -129 237 -123
rect -9 -273 -3 -267
rect -9 -285 -3 -279
rect -9 -297 -3 -291
rect 63 -273 69 -267
rect 63 -285 69 -279
rect 63 -297 69 -291
<< psubdiff >>
rect -60 117 288 120
rect -60 111 -57 117
rect -51 111 -45 117
rect -39 111 -33 117
rect -27 111 -21 117
rect -15 111 -9 117
rect -3 111 3 117
rect 9 111 15 117
rect 21 111 27 117
rect 33 111 39 117
rect 45 111 51 117
rect 57 111 63 117
rect 69 111 75 117
rect 81 111 87 117
rect 93 111 99 117
rect 105 111 111 117
rect 117 111 123 117
rect 129 111 135 117
rect 141 111 147 117
rect 153 111 159 117
rect 165 111 171 117
rect 177 111 183 117
rect 189 111 195 117
rect 201 111 207 117
rect 213 111 219 117
rect 225 111 231 117
rect 237 111 243 117
rect 249 111 255 117
rect 261 111 267 117
rect 273 111 279 117
rect 285 111 288 117
rect -60 108 288 111
rect -60 105 -48 108
rect -60 99 -57 105
rect -51 99 -48 105
rect -60 93 -48 99
rect 108 105 120 108
rect 108 99 111 105
rect 117 99 120 105
rect -60 87 -57 93
rect -51 87 -48 93
rect -60 81 -48 87
rect -60 75 -57 81
rect -51 75 -48 81
rect -60 69 -48 75
rect -60 63 -57 69
rect -51 63 -48 69
rect -60 57 -48 63
rect -60 51 -57 57
rect -51 51 -48 57
rect -60 45 -48 51
rect -60 39 -57 45
rect -51 39 -48 45
rect -60 33 -48 39
rect -60 27 -57 33
rect -51 27 -48 33
rect -60 21 -48 27
rect -60 15 -57 21
rect -51 15 -48 21
rect -60 9 -48 15
rect -60 3 -57 9
rect -51 3 -48 9
rect -60 -3 -48 3
rect -60 -9 -57 -3
rect -51 -9 -48 -3
rect -60 -15 -48 -9
rect -60 -21 -57 -15
rect -51 -21 -48 -15
rect -60 -27 -48 -21
rect 108 93 120 99
rect 276 105 288 108
rect 276 99 279 105
rect 285 99 288 105
rect 108 87 111 93
rect 117 87 120 93
rect 108 81 120 87
rect 108 75 111 81
rect 117 75 120 81
rect 108 69 120 75
rect 108 63 111 69
rect 117 63 120 69
rect 108 57 120 63
rect 108 51 111 57
rect 117 51 120 57
rect 108 45 120 51
rect 108 39 111 45
rect 117 39 120 45
rect 108 33 120 39
rect 108 27 111 33
rect 117 27 120 33
rect 108 21 120 27
rect 108 15 111 21
rect 117 15 120 21
rect 108 9 120 15
rect 108 3 111 9
rect 117 3 120 9
rect 108 -3 120 3
rect 108 -9 111 -3
rect 117 -9 120 -3
rect 108 -15 120 -9
rect 108 -21 111 -15
rect 117 -21 120 -15
rect -60 -33 -57 -27
rect -51 -33 -48 -27
rect -60 -36 -48 -33
rect 108 -27 120 -21
rect 276 93 288 99
rect 276 87 279 93
rect 285 87 288 93
rect 276 81 288 87
rect 276 75 279 81
rect 285 75 288 81
rect 276 69 288 75
rect 276 63 279 69
rect 285 63 288 69
rect 276 57 288 63
rect 276 51 279 57
rect 285 51 288 57
rect 276 45 288 51
rect 276 39 279 45
rect 285 39 288 45
rect 276 33 288 39
rect 276 27 279 33
rect 285 27 288 33
rect 276 21 288 27
rect 276 15 279 21
rect 285 15 288 21
rect 276 9 288 15
rect 276 3 279 9
rect 285 3 288 9
rect 276 -3 288 3
rect 276 -9 279 -3
rect 285 -9 288 -3
rect 276 -15 288 -9
rect 276 -21 279 -15
rect 285 -21 288 -15
rect 108 -33 111 -27
rect 117 -33 120 -27
rect 108 -36 120 -33
rect 276 -27 288 -21
rect 276 -33 279 -27
rect 285 -33 288 -27
rect 276 -36 288 -33
rect -60 -39 288 -36
rect -60 -45 -57 -39
rect -51 -45 -45 -39
rect -39 -45 -33 -39
rect -27 -45 -21 -39
rect -15 -45 -9 -39
rect -3 -45 3 -39
rect 9 -45 15 -39
rect 21 -45 27 -39
rect 33 -45 39 -39
rect 45 -45 51 -39
rect 57 -45 63 -39
rect 69 -45 75 -39
rect 81 -45 87 -39
rect 93 -45 99 -39
rect 105 -45 111 -39
rect 117 -45 123 -39
rect 129 -45 135 -39
rect 141 -45 147 -39
rect 153 -45 159 -39
rect 165 -45 171 -39
rect 177 -45 183 -39
rect 189 -45 195 -39
rect 201 -45 207 -39
rect 213 -45 219 -39
rect 225 -45 231 -39
rect 237 -45 243 -39
rect 249 -45 255 -39
rect 261 -45 267 -39
rect 273 -45 279 -39
rect 285 -45 288 -39
rect -60 -48 288 -45
rect -60 -51 -48 -48
rect -60 -57 -57 -51
rect -51 -57 -48 -51
rect -60 -63 -48 -57
rect 108 -51 120 -48
rect 108 -57 111 -51
rect 117 -57 120 -51
rect -60 -69 -57 -63
rect -51 -69 -48 -63
rect -60 -75 -48 -69
rect -60 -81 -57 -75
rect -51 -81 -48 -75
rect -60 -87 -48 -81
rect -60 -93 -57 -87
rect -51 -93 -48 -87
rect -60 -99 -48 -93
rect -60 -105 -57 -99
rect -51 -105 -48 -99
rect -60 -111 -48 -105
rect -60 -117 -57 -111
rect -51 -117 -48 -111
rect -60 -123 -48 -117
rect -60 -129 -57 -123
rect -51 -129 -48 -123
rect -60 -135 -48 -129
rect -60 -141 -57 -135
rect -51 -141 -48 -135
rect -60 -147 -48 -141
rect -60 -153 -57 -147
rect -51 -153 -48 -147
rect -60 -159 -48 -153
rect -60 -165 -57 -159
rect -51 -165 -48 -159
rect -60 -171 -48 -165
rect -60 -177 -57 -171
rect -51 -177 -48 -171
rect -60 -183 -48 -177
rect 108 -63 120 -57
rect 276 -51 288 -48
rect 276 -57 279 -51
rect 285 -57 288 -51
rect 108 -69 111 -63
rect 117 -69 120 -63
rect 108 -75 120 -69
rect 108 -81 111 -75
rect 117 -81 120 -75
rect 108 -87 120 -81
rect 108 -93 111 -87
rect 117 -93 120 -87
rect 108 -99 120 -93
rect 108 -105 111 -99
rect 117 -105 120 -99
rect 108 -111 120 -105
rect 108 -117 111 -111
rect 117 -117 120 -111
rect 108 -123 120 -117
rect 108 -129 111 -123
rect 117 -129 120 -123
rect 108 -135 120 -129
rect 108 -141 111 -135
rect 117 -141 120 -135
rect 108 -147 120 -141
rect 108 -153 111 -147
rect 117 -153 120 -147
rect 108 -159 120 -153
rect 108 -165 111 -159
rect 117 -165 120 -159
rect 108 -171 120 -165
rect 108 -177 111 -171
rect 117 -177 120 -171
rect -60 -189 -57 -183
rect -51 -189 -48 -183
rect -60 -192 -48 -189
rect 108 -183 120 -177
rect 276 -63 288 -57
rect 276 -69 279 -63
rect 285 -69 288 -63
rect 276 -75 288 -69
rect 276 -81 279 -75
rect 285 -81 288 -75
rect 276 -87 288 -81
rect 276 -93 279 -87
rect 285 -93 288 -87
rect 276 -99 288 -93
rect 276 -105 279 -99
rect 285 -105 288 -99
rect 276 -111 288 -105
rect 276 -117 279 -111
rect 285 -117 288 -111
rect 276 -123 288 -117
rect 276 -129 279 -123
rect 285 -129 288 -123
rect 276 -135 288 -129
rect 276 -141 279 -135
rect 285 -141 288 -135
rect 276 -147 288 -141
rect 276 -153 279 -147
rect 285 -153 288 -147
rect 276 -159 288 -153
rect 276 -165 279 -159
rect 285 -165 288 -159
rect 276 -171 288 -165
rect 276 -177 279 -171
rect 285 -177 288 -171
rect 108 -189 111 -183
rect 117 -189 120 -183
rect 108 -192 120 -189
rect 276 -183 288 -177
rect 276 -189 279 -183
rect 285 -189 288 -183
rect 276 -192 288 -189
rect -60 -195 288 -192
rect -60 -201 -57 -195
rect -51 -201 -45 -195
rect -39 -201 -33 -195
rect -27 -201 -21 -195
rect -15 -201 -9 -195
rect -3 -201 3 -195
rect 9 -201 15 -195
rect 21 -201 27 -195
rect 33 -201 39 -195
rect 45 -201 51 -195
rect 57 -201 63 -195
rect 69 -201 75 -195
rect 81 -201 87 -195
rect 93 -201 99 -195
rect 105 -201 111 -195
rect 117 -201 123 -195
rect 129 -201 135 -195
rect 141 -201 147 -195
rect 153 -201 159 -195
rect 165 -201 171 -195
rect 177 -201 183 -195
rect 189 -201 195 -195
rect 201 -201 207 -195
rect 213 -201 219 -195
rect 225 -201 231 -195
rect 237 -201 243 -195
rect 249 -201 255 -195
rect 261 -201 267 -195
rect 273 -201 279 -195
rect 285 -201 288 -195
rect -60 -204 288 -201
rect -60 -207 -48 -204
rect -60 -213 -57 -207
rect -51 -213 -48 -207
rect -60 -219 -48 -213
rect 108 -207 120 -204
rect 108 -213 111 -207
rect 117 -213 120 -207
rect -60 -225 -57 -219
rect -51 -225 -48 -219
rect -60 -231 -48 -225
rect -60 -237 -57 -231
rect -51 -237 -48 -231
rect -60 -243 -48 -237
rect -60 -249 -57 -243
rect -51 -249 -48 -243
rect -60 -255 -48 -249
rect -60 -261 -57 -255
rect -51 -261 -48 -255
rect -60 -267 -48 -261
rect -60 -273 -57 -267
rect -51 -273 -48 -267
rect -60 -279 -48 -273
rect -60 -285 -57 -279
rect -51 -285 -48 -279
rect -60 -291 -48 -285
rect -60 -297 -57 -291
rect -51 -297 -48 -291
rect -60 -303 -48 -297
rect -60 -309 -57 -303
rect -51 -309 -48 -303
rect -60 -315 -48 -309
rect -60 -321 -57 -315
rect -51 -321 -48 -315
rect -60 -327 -48 -321
rect -60 -333 -57 -327
rect -51 -333 -48 -327
rect -60 -339 -48 -333
rect 108 -219 120 -213
rect 108 -225 111 -219
rect 117 -225 120 -219
rect 108 -231 120 -225
rect 108 -237 111 -231
rect 117 -237 120 -231
rect 108 -243 120 -237
rect 276 -207 288 -204
rect 276 -213 279 -207
rect 285 -213 288 -207
rect 276 -219 288 -213
rect 276 -225 279 -219
rect 285 -225 288 -219
rect 276 -231 288 -225
rect 276 -237 279 -231
rect 285 -237 288 -231
rect 108 -249 111 -243
rect 117 -249 120 -243
rect 108 -255 120 -249
rect 108 -261 111 -255
rect 117 -261 120 -255
rect 108 -267 120 -261
rect 276 -243 288 -237
rect 276 -249 279 -243
rect 285 -249 288 -243
rect 276 -255 288 -249
rect 276 -261 279 -255
rect 285 -261 288 -255
rect 108 -273 111 -267
rect 117 -273 120 -267
rect 108 -279 120 -273
rect 108 -285 111 -279
rect 117 -285 120 -279
rect 108 -291 120 -285
rect 108 -297 111 -291
rect 117 -297 120 -291
rect 108 -303 120 -297
rect 276 -267 288 -261
rect 276 -273 279 -267
rect 285 -273 288 -267
rect 276 -279 288 -273
rect 276 -285 279 -279
rect 285 -285 288 -279
rect 276 -291 288 -285
rect 276 -297 279 -291
rect 285 -297 288 -291
rect 108 -309 111 -303
rect 117 -309 120 -303
rect 276 -303 288 -297
rect 108 -315 120 -309
rect 108 -321 111 -315
rect 117 -321 120 -315
rect 108 -327 120 -321
rect 108 -333 111 -327
rect 117 -333 120 -327
rect -60 -345 -57 -339
rect -51 -345 -48 -339
rect -60 -348 -48 -345
rect 108 -339 120 -333
rect 108 -345 111 -339
rect 117 -345 120 -339
rect 108 -348 120 -345
rect 276 -309 279 -303
rect 285 -309 288 -303
rect 276 -315 288 -309
rect 276 -321 279 -315
rect 285 -321 288 -315
rect 276 -327 288 -321
rect 276 -333 279 -327
rect 285 -333 288 -327
rect 276 -339 288 -333
rect 276 -345 279 -339
rect 285 -345 288 -339
rect 276 -348 288 -345
rect -60 -351 288 -348
rect -60 -357 -57 -351
rect -51 -357 -45 -351
rect -39 -357 -33 -351
rect -27 -357 -21 -351
rect -15 -357 -9 -351
rect -3 -357 3 -351
rect 9 -357 15 -351
rect 21 -357 27 -351
rect 33 -357 39 -351
rect 45 -357 51 -351
rect 57 -357 63 -351
rect 69 -357 75 -351
rect 81 -357 87 -351
rect 93 -357 99 -351
rect 105 -357 111 -351
rect 117 -357 123 -351
rect 129 -357 135 -351
rect 141 -357 147 -351
rect 153 -357 159 -351
rect 165 -357 171 -351
rect 177 -357 183 -351
rect 189 -357 195 -351
rect 201 -357 207 -351
rect 213 -357 219 -351
rect 225 -357 231 -351
rect 237 -357 243 -351
rect 249 -357 255 -351
rect 261 -357 267 -351
rect 273 -357 279 -351
rect 285 -357 288 -351
rect -60 -360 288 -357
<< nsubdiff >>
rect -36 93 96 96
rect -36 87 -33 93
rect -27 87 -21 93
rect -15 87 -9 93
rect -3 87 3 93
rect 9 87 15 93
rect 21 87 27 93
rect 33 87 39 93
rect 45 87 51 93
rect 57 87 63 93
rect 69 87 75 93
rect 81 87 87 93
rect 93 87 96 93
rect -36 84 96 87
rect -36 81 -24 84
rect -36 75 -33 81
rect -27 75 -24 81
rect -36 69 -24 75
rect 84 81 96 84
rect 84 75 87 81
rect 93 75 96 81
rect -36 63 -33 69
rect -27 63 -24 69
rect -36 57 -24 63
rect -36 51 -33 57
rect -27 51 -24 57
rect -36 45 -24 51
rect 84 69 96 75
rect 84 63 87 69
rect 93 63 96 69
rect 84 57 96 63
rect 84 51 87 57
rect 93 51 96 57
rect -36 39 -33 45
rect -27 39 -24 45
rect -36 33 -24 39
rect -36 27 -33 33
rect -27 27 -24 33
rect -36 21 -24 27
rect -36 15 -33 21
rect -27 15 -24 21
rect -36 9 -24 15
rect 84 45 96 51
rect 84 39 87 45
rect 93 39 96 45
rect 84 33 96 39
rect 84 27 87 33
rect 93 27 96 33
rect 84 21 96 27
rect 84 15 87 21
rect 93 15 96 21
rect -36 3 -33 9
rect -27 3 -24 9
rect 84 9 96 15
rect -36 -3 -24 3
rect -36 -9 -33 -3
rect -27 -9 -24 -3
rect -36 -12 -24 -9
rect 84 3 87 9
rect 93 3 96 9
rect 84 -3 96 3
rect 84 -9 87 -3
rect 93 -9 96 -3
rect 84 -12 96 -9
rect -36 -15 96 -12
rect -36 -21 -33 -15
rect -27 -21 -21 -15
rect -15 -21 -9 -15
rect -3 -21 3 -15
rect 9 -21 15 -15
rect 21 -21 27 -15
rect 33 -21 39 -15
rect 45 -21 51 -15
rect 57 -21 63 -15
rect 69 -21 75 -15
rect 81 -21 87 -15
rect 93 -21 96 -15
rect -36 -24 96 -21
rect 132 93 264 96
rect 132 87 135 93
rect 141 87 147 93
rect 153 87 159 93
rect 165 87 171 93
rect 177 87 183 93
rect 189 87 195 93
rect 201 87 207 93
rect 213 87 219 93
rect 225 87 231 93
rect 237 87 243 93
rect 249 87 255 93
rect 261 87 264 93
rect 132 84 264 87
rect 132 81 144 84
rect 132 75 135 81
rect 141 75 144 81
rect 132 69 144 75
rect 252 81 264 84
rect 252 75 255 81
rect 261 75 264 81
rect 132 63 135 69
rect 141 63 144 69
rect 132 57 144 63
rect 132 51 135 57
rect 141 51 144 57
rect 132 45 144 51
rect 252 69 264 75
rect 252 63 255 69
rect 261 63 264 69
rect 252 57 264 63
rect 252 51 255 57
rect 261 51 264 57
rect 132 39 135 45
rect 141 39 144 45
rect 132 33 144 39
rect 132 27 135 33
rect 141 27 144 33
rect 132 21 144 27
rect 132 15 135 21
rect 141 15 144 21
rect 132 9 144 15
rect 252 45 264 51
rect 252 39 255 45
rect 261 39 264 45
rect 252 33 264 39
rect 252 27 255 33
rect 261 27 264 33
rect 252 21 264 27
rect 252 15 255 21
rect 261 15 264 21
rect 132 3 135 9
rect 141 3 144 9
rect 252 9 264 15
rect 132 -3 144 3
rect 132 -9 135 -3
rect 141 -9 144 -3
rect 132 -12 144 -9
rect 252 3 255 9
rect 261 3 264 9
rect 252 -3 264 3
rect 252 -9 255 -3
rect 261 -9 264 -3
rect 252 -12 264 -9
rect 132 -15 264 -12
rect 132 -21 135 -15
rect 141 -21 147 -15
rect 153 -21 159 -15
rect 165 -21 171 -15
rect 177 -21 183 -15
rect 189 -21 195 -15
rect 201 -21 207 -15
rect 213 -21 219 -15
rect 225 -21 231 -15
rect 237 -21 243 -15
rect 249 -21 255 -15
rect 261 -21 264 -15
rect 132 -24 264 -21
rect -36 -63 96 -60
rect -36 -69 -33 -63
rect -27 -69 -21 -63
rect -15 -69 -9 -63
rect -3 -69 3 -63
rect 9 -69 15 -63
rect 21 -69 27 -63
rect 33 -69 39 -63
rect 45 -69 51 -63
rect 57 -69 63 -63
rect 69 -69 75 -63
rect 81 -69 87 -63
rect 93 -69 96 -63
rect -36 -72 96 -69
rect -36 -75 -24 -72
rect -36 -81 -33 -75
rect -27 -81 -24 -75
rect -36 -87 -24 -81
rect -36 -93 -33 -87
rect -27 -93 -24 -87
rect 84 -75 96 -72
rect 84 -81 87 -75
rect 93 -81 96 -75
rect 84 -87 96 -81
rect -36 -99 -24 -93
rect 84 -93 87 -87
rect 93 -93 96 -87
rect -36 -105 -33 -99
rect -27 -105 -24 -99
rect -36 -111 -24 -105
rect -36 -117 -33 -111
rect -27 -117 -24 -111
rect -36 -123 -24 -117
rect -36 -129 -33 -123
rect -27 -129 -24 -123
rect -36 -135 -24 -129
rect 84 -99 96 -93
rect 84 -105 87 -99
rect 93 -105 96 -99
rect 84 -111 96 -105
rect 84 -117 87 -111
rect 93 -117 96 -111
rect 84 -123 96 -117
rect 84 -129 87 -123
rect 93 -129 96 -123
rect -36 -141 -33 -135
rect -27 -141 -24 -135
rect -36 -147 -24 -141
rect -36 -153 -33 -147
rect -27 -153 -24 -147
rect -36 -159 -24 -153
rect 84 -135 96 -129
rect 84 -141 87 -135
rect 93 -141 96 -135
rect 84 -147 96 -141
rect 84 -153 87 -147
rect 93 -153 96 -147
rect -36 -165 -33 -159
rect -27 -165 -24 -159
rect -36 -168 -24 -165
rect 84 -159 96 -153
rect 84 -165 87 -159
rect 93 -165 96 -159
rect 84 -168 96 -165
rect -36 -171 96 -168
rect -36 -177 -33 -171
rect -27 -177 -21 -171
rect -15 -177 -9 -171
rect -3 -177 3 -171
rect 9 -177 15 -171
rect 21 -177 27 -171
rect 33 -177 39 -171
rect 45 -177 51 -171
rect 57 -177 63 -171
rect 69 -177 75 -171
rect 81 -177 87 -171
rect 93 -177 96 -171
rect -36 -180 96 -177
rect 132 -63 264 -60
rect 132 -69 135 -63
rect 141 -69 147 -63
rect 153 -69 159 -63
rect 165 -69 171 -63
rect 177 -69 183 -63
rect 189 -69 195 -63
rect 201 -69 207 -63
rect 213 -69 219 -63
rect 225 -69 231 -63
rect 237 -69 243 -63
rect 249 -69 255 -63
rect 261 -69 264 -63
rect 132 -72 264 -69
rect 132 -75 144 -72
rect 132 -81 135 -75
rect 141 -81 144 -75
rect 132 -87 144 -81
rect 132 -93 135 -87
rect 141 -93 144 -87
rect 252 -75 264 -72
rect 252 -81 255 -75
rect 261 -81 264 -75
rect 252 -87 264 -81
rect 132 -99 144 -93
rect 252 -93 255 -87
rect 261 -93 264 -87
rect 132 -105 135 -99
rect 141 -105 144 -99
rect 132 -111 144 -105
rect 132 -117 135 -111
rect 141 -117 144 -111
rect 132 -123 144 -117
rect 132 -129 135 -123
rect 141 -129 144 -123
rect 132 -135 144 -129
rect 252 -99 264 -93
rect 252 -105 255 -99
rect 261 -105 264 -99
rect 252 -111 264 -105
rect 252 -117 255 -111
rect 261 -117 264 -111
rect 252 -123 264 -117
rect 252 -129 255 -123
rect 261 -129 264 -123
rect 132 -141 135 -135
rect 141 -141 144 -135
rect 132 -147 144 -141
rect 132 -153 135 -147
rect 141 -153 144 -147
rect 132 -159 144 -153
rect 252 -135 264 -129
rect 252 -141 255 -135
rect 261 -141 264 -135
rect 252 -147 264 -141
rect 252 -153 255 -147
rect 261 -153 264 -147
rect 132 -165 135 -159
rect 141 -165 144 -159
rect 132 -168 144 -165
rect 252 -159 264 -153
rect 252 -165 255 -159
rect 261 -165 264 -159
rect 252 -168 264 -165
rect 132 -171 264 -168
rect 132 -177 135 -171
rect 141 -177 147 -171
rect 153 -177 159 -171
rect 165 -177 171 -171
rect 177 -177 183 -171
rect 189 -177 195 -171
rect 201 -177 207 -171
rect 213 -177 219 -171
rect 225 -177 231 -171
rect 237 -177 243 -171
rect 249 -177 255 -171
rect 261 -177 264 -171
rect 132 -180 264 -177
rect -36 -219 96 -216
rect -36 -225 -33 -219
rect -27 -225 -21 -219
rect -15 -225 -9 -219
rect -3 -225 3 -219
rect 9 -225 15 -219
rect 21 -225 27 -219
rect 33 -225 39 -219
rect 45 -225 51 -219
rect 57 -225 63 -219
rect 69 -225 75 -219
rect 81 -225 87 -219
rect 93 -225 96 -219
rect -36 -228 96 -225
rect -36 -231 -24 -228
rect -36 -237 -33 -231
rect -27 -237 -24 -231
rect -36 -243 -24 -237
rect 84 -231 96 -228
rect 84 -237 87 -231
rect 93 -237 96 -231
rect -36 -249 -33 -243
rect -27 -249 -24 -243
rect -36 -255 -24 -249
rect -36 -261 -33 -255
rect -27 -261 -24 -255
rect -36 -267 -24 -261
rect 84 -243 96 -237
rect 84 -249 87 -243
rect 93 -249 96 -243
rect 84 -255 96 -249
rect 84 -261 87 -255
rect 93 -261 96 -255
rect -36 -273 -33 -267
rect -27 -273 -24 -267
rect -36 -279 -24 -273
rect -36 -285 -33 -279
rect -27 -285 -24 -279
rect -36 -291 -24 -285
rect -36 -297 -33 -291
rect -27 -297 -24 -291
rect -36 -303 -24 -297
rect 84 -267 96 -261
rect 84 -273 87 -267
rect 93 -273 96 -267
rect 84 -279 96 -273
rect 84 -285 87 -279
rect 93 -285 96 -279
rect 84 -291 96 -285
rect 84 -297 87 -291
rect 93 -297 96 -291
rect -36 -309 -33 -303
rect -27 -309 -24 -303
rect 84 -303 96 -297
rect -36 -315 -24 -309
rect -36 -321 -33 -315
rect -27 -321 -24 -315
rect -36 -324 -24 -321
rect 84 -309 87 -303
rect 93 -309 96 -303
rect 84 -315 96 -309
rect 84 -321 87 -315
rect 93 -321 96 -315
rect 84 -324 96 -321
rect -36 -327 96 -324
rect -36 -333 -33 -327
rect -27 -333 -21 -327
rect -15 -333 -9 -327
rect -3 -333 3 -327
rect 9 -333 15 -327
rect 21 -333 27 -327
rect 33 -333 39 -327
rect 45 -333 51 -327
rect 57 -333 63 -327
rect 69 -333 75 -327
rect 81 -333 87 -327
rect 93 -333 96 -327
rect -36 -336 96 -333
<< psubdiffcont >>
rect -57 111 -51 117
rect -45 111 -39 117
rect -33 111 -27 117
rect -21 111 -15 117
rect -9 111 -3 117
rect 3 111 9 117
rect 15 111 21 117
rect 27 111 33 117
rect 39 111 45 117
rect 51 111 57 117
rect 63 111 69 117
rect 75 111 81 117
rect 87 111 93 117
rect 99 111 105 117
rect 111 111 117 117
rect 123 111 129 117
rect 135 111 141 117
rect 147 111 153 117
rect 159 111 165 117
rect 171 111 177 117
rect 183 111 189 117
rect 195 111 201 117
rect 207 111 213 117
rect 219 111 225 117
rect 231 111 237 117
rect 243 111 249 117
rect 255 111 261 117
rect 267 111 273 117
rect 279 111 285 117
rect -57 99 -51 105
rect 111 99 117 105
rect -57 87 -51 93
rect -57 75 -51 81
rect -57 63 -51 69
rect -57 51 -51 57
rect -57 39 -51 45
rect -57 27 -51 33
rect -57 15 -51 21
rect -57 3 -51 9
rect -57 -9 -51 -3
rect -57 -21 -51 -15
rect 279 99 285 105
rect 111 87 117 93
rect 111 75 117 81
rect 111 63 117 69
rect 111 51 117 57
rect 111 39 117 45
rect 111 27 117 33
rect 111 15 117 21
rect 111 3 117 9
rect 111 -9 117 -3
rect 111 -21 117 -15
rect -57 -33 -51 -27
rect 279 87 285 93
rect 279 75 285 81
rect 279 63 285 69
rect 279 51 285 57
rect 279 39 285 45
rect 279 27 285 33
rect 279 15 285 21
rect 279 3 285 9
rect 279 -9 285 -3
rect 279 -21 285 -15
rect 111 -33 117 -27
rect 279 -33 285 -27
rect -57 -45 -51 -39
rect -45 -45 -39 -39
rect -33 -45 -27 -39
rect -21 -45 -15 -39
rect -9 -45 -3 -39
rect 3 -45 9 -39
rect 15 -45 21 -39
rect 27 -45 33 -39
rect 39 -45 45 -39
rect 51 -45 57 -39
rect 63 -45 69 -39
rect 75 -45 81 -39
rect 87 -45 93 -39
rect 99 -45 105 -39
rect 111 -45 117 -39
rect 123 -45 129 -39
rect 135 -45 141 -39
rect 147 -45 153 -39
rect 159 -45 165 -39
rect 171 -45 177 -39
rect 183 -45 189 -39
rect 195 -45 201 -39
rect 207 -45 213 -39
rect 219 -45 225 -39
rect 231 -45 237 -39
rect 243 -45 249 -39
rect 255 -45 261 -39
rect 267 -45 273 -39
rect 279 -45 285 -39
rect -57 -57 -51 -51
rect 111 -57 117 -51
rect -57 -69 -51 -63
rect -57 -81 -51 -75
rect -57 -93 -51 -87
rect -57 -105 -51 -99
rect -57 -117 -51 -111
rect -57 -129 -51 -123
rect -57 -141 -51 -135
rect -57 -153 -51 -147
rect -57 -165 -51 -159
rect -57 -177 -51 -171
rect 279 -57 285 -51
rect 111 -69 117 -63
rect 111 -81 117 -75
rect 111 -93 117 -87
rect 111 -105 117 -99
rect 111 -117 117 -111
rect 111 -129 117 -123
rect 111 -141 117 -135
rect 111 -153 117 -147
rect 111 -165 117 -159
rect 111 -177 117 -171
rect -57 -189 -51 -183
rect 279 -69 285 -63
rect 279 -81 285 -75
rect 279 -93 285 -87
rect 279 -105 285 -99
rect 279 -117 285 -111
rect 279 -129 285 -123
rect 279 -141 285 -135
rect 279 -153 285 -147
rect 279 -165 285 -159
rect 279 -177 285 -171
rect 111 -189 117 -183
rect 279 -189 285 -183
rect -57 -201 -51 -195
rect -45 -201 -39 -195
rect -33 -201 -27 -195
rect -21 -201 -15 -195
rect -9 -201 -3 -195
rect 3 -201 9 -195
rect 15 -201 21 -195
rect 27 -201 33 -195
rect 39 -201 45 -195
rect 51 -201 57 -195
rect 63 -201 69 -195
rect 75 -201 81 -195
rect 87 -201 93 -195
rect 99 -201 105 -195
rect 111 -201 117 -195
rect 123 -201 129 -195
rect 135 -201 141 -195
rect 147 -201 153 -195
rect 159 -201 165 -195
rect 171 -201 177 -195
rect 183 -201 189 -195
rect 195 -201 201 -195
rect 207 -201 213 -195
rect 219 -201 225 -195
rect 231 -201 237 -195
rect 243 -201 249 -195
rect 255 -201 261 -195
rect 267 -201 273 -195
rect 279 -201 285 -195
rect -57 -213 -51 -207
rect 111 -213 117 -207
rect -57 -225 -51 -219
rect -57 -237 -51 -231
rect -57 -249 -51 -243
rect -57 -261 -51 -255
rect -57 -273 -51 -267
rect -57 -285 -51 -279
rect -57 -297 -51 -291
rect -57 -309 -51 -303
rect -57 -321 -51 -315
rect -57 -333 -51 -327
rect 111 -225 117 -219
rect 111 -237 117 -231
rect 279 -213 285 -207
rect 279 -225 285 -219
rect 279 -237 285 -231
rect 111 -249 117 -243
rect 111 -261 117 -255
rect 279 -249 285 -243
rect 279 -261 285 -255
rect 111 -273 117 -267
rect 111 -285 117 -279
rect 111 -297 117 -291
rect 279 -273 285 -267
rect 279 -285 285 -279
rect 279 -297 285 -291
rect 111 -309 117 -303
rect 111 -321 117 -315
rect 111 -333 117 -327
rect -57 -345 -51 -339
rect 111 -345 117 -339
rect 279 -309 285 -303
rect 279 -321 285 -315
rect 279 -333 285 -327
rect 279 -345 285 -339
rect -57 -357 -51 -351
rect -45 -357 -39 -351
rect -33 -357 -27 -351
rect -21 -357 -15 -351
rect -9 -357 -3 -351
rect 3 -357 9 -351
rect 15 -357 21 -351
rect 27 -357 33 -351
rect 39 -357 45 -351
rect 51 -357 57 -351
rect 63 -357 69 -351
rect 75 -357 81 -351
rect 87 -357 93 -351
rect 99 -357 105 -351
rect 111 -357 117 -351
rect 123 -357 129 -351
rect 135 -357 141 -351
rect 147 -357 153 -351
rect 159 -357 165 -351
rect 171 -357 177 -351
rect 183 -357 189 -351
rect 195 -357 201 -351
rect 207 -357 213 -351
rect 219 -357 225 -351
rect 231 -357 237 -351
rect 243 -357 249 -351
rect 255 -357 261 -351
rect 267 -357 273 -351
rect 279 -357 285 -351
<< nsubdiffcont >>
rect -33 87 -27 93
rect -21 87 -15 93
rect -9 87 -3 93
rect 3 87 9 93
rect 15 87 21 93
rect 27 87 33 93
rect 39 87 45 93
rect 51 87 57 93
rect 63 87 69 93
rect 75 87 81 93
rect 87 87 93 93
rect -33 75 -27 81
rect 87 75 93 81
rect -33 63 -27 69
rect -33 51 -27 57
rect 87 63 93 69
rect 87 51 93 57
rect -33 39 -27 45
rect -33 27 -27 33
rect -33 15 -27 21
rect 87 39 93 45
rect 87 27 93 33
rect 87 15 93 21
rect -33 3 -27 9
rect -33 -9 -27 -3
rect 87 3 93 9
rect 87 -9 93 -3
rect -33 -21 -27 -15
rect -21 -21 -15 -15
rect -9 -21 -3 -15
rect 3 -21 9 -15
rect 15 -21 21 -15
rect 27 -21 33 -15
rect 39 -21 45 -15
rect 51 -21 57 -15
rect 63 -21 69 -15
rect 75 -21 81 -15
rect 87 -21 93 -15
rect 135 87 141 93
rect 147 87 153 93
rect 159 87 165 93
rect 171 87 177 93
rect 183 87 189 93
rect 195 87 201 93
rect 207 87 213 93
rect 219 87 225 93
rect 231 87 237 93
rect 243 87 249 93
rect 255 87 261 93
rect 135 75 141 81
rect 255 75 261 81
rect 135 63 141 69
rect 135 51 141 57
rect 255 63 261 69
rect 255 51 261 57
rect 135 39 141 45
rect 135 27 141 33
rect 135 15 141 21
rect 255 39 261 45
rect 255 27 261 33
rect 255 15 261 21
rect 135 3 141 9
rect 135 -9 141 -3
rect 255 3 261 9
rect 255 -9 261 -3
rect 135 -21 141 -15
rect 147 -21 153 -15
rect 159 -21 165 -15
rect 171 -21 177 -15
rect 183 -21 189 -15
rect 195 -21 201 -15
rect 207 -21 213 -15
rect 219 -21 225 -15
rect 231 -21 237 -15
rect 243 -21 249 -15
rect 255 -21 261 -15
rect -33 -69 -27 -63
rect -21 -69 -15 -63
rect -9 -69 -3 -63
rect 3 -69 9 -63
rect 15 -69 21 -63
rect 27 -69 33 -63
rect 39 -69 45 -63
rect 51 -69 57 -63
rect 63 -69 69 -63
rect 75 -69 81 -63
rect 87 -69 93 -63
rect -33 -81 -27 -75
rect -33 -93 -27 -87
rect 87 -81 93 -75
rect 87 -93 93 -87
rect -33 -105 -27 -99
rect -33 -117 -27 -111
rect -33 -129 -27 -123
rect 87 -105 93 -99
rect 87 -117 93 -111
rect 87 -129 93 -123
rect -33 -141 -27 -135
rect -33 -153 -27 -147
rect 87 -141 93 -135
rect 87 -153 93 -147
rect -33 -165 -27 -159
rect 87 -165 93 -159
rect -33 -177 -27 -171
rect -21 -177 -15 -171
rect -9 -177 -3 -171
rect 3 -177 9 -171
rect 15 -177 21 -171
rect 27 -177 33 -171
rect 39 -177 45 -171
rect 51 -177 57 -171
rect 63 -177 69 -171
rect 75 -177 81 -171
rect 87 -177 93 -171
rect 135 -69 141 -63
rect 147 -69 153 -63
rect 159 -69 165 -63
rect 171 -69 177 -63
rect 183 -69 189 -63
rect 195 -69 201 -63
rect 207 -69 213 -63
rect 219 -69 225 -63
rect 231 -69 237 -63
rect 243 -69 249 -63
rect 255 -69 261 -63
rect 135 -81 141 -75
rect 135 -93 141 -87
rect 255 -81 261 -75
rect 255 -93 261 -87
rect 135 -105 141 -99
rect 135 -117 141 -111
rect 135 -129 141 -123
rect 255 -105 261 -99
rect 255 -117 261 -111
rect 255 -129 261 -123
rect 135 -141 141 -135
rect 135 -153 141 -147
rect 255 -141 261 -135
rect 255 -153 261 -147
rect 135 -165 141 -159
rect 255 -165 261 -159
rect 135 -177 141 -171
rect 147 -177 153 -171
rect 159 -177 165 -171
rect 171 -177 177 -171
rect 183 -177 189 -171
rect 195 -177 201 -171
rect 207 -177 213 -171
rect 219 -177 225 -171
rect 231 -177 237 -171
rect 243 -177 249 -171
rect 255 -177 261 -171
rect -33 -225 -27 -219
rect -21 -225 -15 -219
rect -9 -225 -3 -219
rect 3 -225 9 -219
rect 15 -225 21 -219
rect 27 -225 33 -219
rect 39 -225 45 -219
rect 51 -225 57 -219
rect 63 -225 69 -219
rect 75 -225 81 -219
rect 87 -225 93 -219
rect -33 -237 -27 -231
rect 87 -237 93 -231
rect -33 -249 -27 -243
rect -33 -261 -27 -255
rect 87 -249 93 -243
rect 87 -261 93 -255
rect -33 -273 -27 -267
rect -33 -285 -27 -279
rect -33 -297 -27 -291
rect 87 -273 93 -267
rect 87 -285 93 -279
rect 87 -297 93 -291
rect -33 -309 -27 -303
rect -33 -321 -27 -315
rect 87 -309 93 -303
rect 87 -321 93 -315
rect -33 -333 -27 -327
rect -21 -333 -15 -327
rect -9 -333 -3 -327
rect 3 -333 9 -327
rect 15 -333 21 -327
rect 27 -333 33 -327
rect 39 -333 45 -327
rect 51 -333 57 -327
rect 63 -333 69 -327
rect 75 -333 81 -327
rect 87 -333 93 -327
<< polysilicon >>
rect 0 69 60 72
rect 0 63 3 69
rect 9 63 15 69
rect 21 63 27 69
rect 33 63 39 69
rect 45 63 51 69
rect 57 63 60 69
rect 0 48 60 63
rect 0 6 60 12
rect 168 69 228 72
rect 168 63 171 69
rect 177 63 183 69
rect 189 63 195 69
rect 201 63 207 69
rect 213 63 219 69
rect 225 63 228 69
rect 168 48 228 63
rect 168 6 228 12
rect 0 -96 60 -90
rect 0 -147 60 -132
rect 0 -153 3 -147
rect 9 -153 15 -147
rect 21 -153 27 -147
rect 33 -153 39 -147
rect 45 -153 51 -147
rect 57 -153 60 -147
rect 0 -156 60 -153
rect 168 -96 228 -90
rect 168 -147 228 -132
rect 168 -153 171 -147
rect 177 -153 183 -147
rect 189 -153 195 -147
rect 201 -153 207 -147
rect 213 -153 219 -147
rect 225 -153 228 -147
rect 168 -156 228 -153
rect 0 -243 60 -240
rect 0 -249 3 -243
rect 9 -249 15 -243
rect 21 -249 27 -243
rect 33 -249 39 -243
rect 45 -249 51 -243
rect 57 -249 60 -243
rect 0 -264 60 -249
rect 0 -306 60 -300
rect 168 -243 228 -240
rect 168 -249 171 -243
rect 177 -249 183 -243
rect 189 -249 195 -243
rect 201 -249 207 -243
rect 213 -249 219 -243
rect 225 -249 228 -243
rect 168 -264 228 -249
rect 168 -306 228 -300
<< polycontact >>
rect 3 63 9 69
rect 15 63 21 69
rect 27 63 33 69
rect 39 63 45 69
rect 51 63 57 69
rect 171 63 177 69
rect 183 63 189 69
rect 195 63 201 69
rect 207 63 213 69
rect 219 63 225 69
rect 3 -153 9 -147
rect 15 -153 21 -147
rect 27 -153 33 -147
rect 39 -153 45 -147
rect 51 -153 57 -147
rect 171 -153 177 -147
rect 183 -153 189 -147
rect 195 -153 201 -147
rect 207 -153 213 -147
rect 219 -153 225 -147
rect 3 -249 9 -243
rect 15 -249 21 -243
rect 27 -249 33 -243
rect 39 -249 45 -243
rect 51 -249 57 -243
rect 171 -249 177 -243
rect 183 -249 189 -243
rect 195 -249 201 -243
rect 207 -249 213 -243
rect 219 -249 225 -243
<< metal1 >>
rect -60 117 288 120
rect -60 111 -57 117
rect -51 111 -45 117
rect -39 111 -33 117
rect -27 111 -21 117
rect -15 111 -9 117
rect -3 111 3 117
rect 9 111 15 117
rect 21 111 27 117
rect 33 111 39 117
rect 45 111 51 117
rect 57 111 63 117
rect 69 111 75 117
rect 81 111 87 117
rect 93 111 99 117
rect 105 111 111 117
rect 117 111 123 117
rect 129 111 135 117
rect 141 111 147 117
rect 153 111 159 117
rect 165 111 171 117
rect 177 111 183 117
rect 189 111 195 117
rect 201 111 207 117
rect 213 111 219 117
rect 225 111 231 117
rect 237 111 243 117
rect 249 111 255 117
rect 261 111 267 117
rect 273 111 279 117
rect 285 111 288 117
rect -60 108 288 111
rect -60 105 -48 108
rect -60 99 -57 105
rect -51 99 -48 105
rect -60 93 -48 99
rect 108 105 120 108
rect 108 99 111 105
rect 117 99 120 105
rect -60 87 -57 93
rect -51 87 -48 93
rect -60 81 -48 87
rect -60 75 -57 81
rect -51 75 -48 81
rect -60 69 -48 75
rect -60 63 -57 69
rect -51 63 -48 69
rect -60 57 -48 63
rect -60 51 -57 57
rect -51 51 -48 57
rect -60 45 -48 51
rect -60 39 -57 45
rect -51 39 -48 45
rect -60 33 -48 39
rect -60 27 -57 33
rect -51 27 -48 33
rect -60 21 -48 27
rect -60 15 -57 21
rect -51 15 -48 21
rect -60 9 -48 15
rect -60 3 -57 9
rect -51 3 -48 9
rect -60 -3 -48 3
rect -60 -9 -57 -3
rect -51 -9 -48 -3
rect -60 -15 -48 -9
rect -60 -21 -57 -15
rect -51 -21 -48 -15
rect -60 -27 -48 -21
rect -36 93 96 96
rect -36 87 -33 93
rect -27 87 -21 93
rect -15 87 -9 93
rect -3 87 3 93
rect 9 87 15 93
rect 21 87 27 93
rect 33 87 39 93
rect 45 87 51 93
rect 57 87 63 93
rect 69 87 75 93
rect 81 87 87 93
rect 93 87 96 93
rect -36 84 96 87
rect -36 81 -24 84
rect -36 75 -33 81
rect -27 75 -24 81
rect -36 69 -24 75
rect 84 81 96 84
rect 84 75 87 81
rect 93 75 96 81
rect -36 63 -33 69
rect -27 63 -24 69
rect -36 57 -24 63
rect -36 51 -33 57
rect -27 51 -24 57
rect -36 45 -24 51
rect -36 39 -33 45
rect -27 39 -24 45
rect -36 33 -24 39
rect -36 27 -33 33
rect -27 27 -24 33
rect -36 21 -24 27
rect -36 15 -33 21
rect -27 15 -24 21
rect -36 9 -24 15
rect -12 69 60 72
rect -12 63 -9 69
rect -3 63 3 69
rect 9 63 15 69
rect 21 63 27 69
rect 33 63 39 69
rect 45 63 51 69
rect 57 63 60 69
rect -12 60 60 63
rect 84 69 96 75
rect 84 63 87 69
rect 93 63 96 69
rect -12 57 0 60
rect -12 51 -9 57
rect -3 51 0 57
rect -12 45 0 51
rect 84 57 96 63
rect 84 51 87 57
rect 93 51 96 57
rect -12 39 -9 45
rect -3 39 0 45
rect -12 33 0 39
rect -12 27 -9 33
rect -3 27 0 33
rect -12 21 0 27
rect -12 15 -9 21
rect -3 15 0 21
rect -12 12 0 15
rect 60 45 72 48
rect 60 39 63 45
rect 69 39 72 45
rect 60 33 72 39
rect 60 27 63 33
rect 69 27 72 33
rect 60 21 72 27
rect 60 15 63 21
rect 69 15 72 21
rect -36 3 -33 9
rect -27 3 -24 9
rect -36 -3 -24 3
rect -36 -9 -33 -3
rect -27 -9 -24 -3
rect -36 -12 -24 -9
rect 60 -12 72 15
rect 84 45 96 51
rect 84 39 87 45
rect 93 39 96 45
rect 84 33 96 39
rect 84 27 87 33
rect 93 27 96 33
rect 84 21 96 27
rect 84 15 87 21
rect 93 15 96 21
rect 84 9 96 15
rect 84 3 87 9
rect 93 3 96 9
rect 84 -3 96 3
rect 84 -9 87 -3
rect 93 -9 96 -3
rect 84 -12 96 -9
rect -36 -15 96 -12
rect -36 -21 -33 -15
rect -27 -21 -21 -15
rect -15 -21 -9 -15
rect -3 -21 3 -15
rect 9 -21 15 -15
rect 21 -21 27 -15
rect 33 -21 39 -15
rect 45 -21 51 -15
rect 57 -21 63 -15
rect 69 -21 75 -15
rect 81 -21 87 -15
rect 93 -21 96 -15
rect -36 -24 96 -21
rect 108 93 120 99
rect 276 105 288 108
rect 276 99 279 105
rect 285 99 288 105
rect 108 87 111 93
rect 117 87 120 93
rect 108 81 120 87
rect 108 75 111 81
rect 117 75 120 81
rect 108 69 120 75
rect 108 63 111 69
rect 117 63 120 69
rect 108 57 120 63
rect 108 51 111 57
rect 117 51 120 57
rect 108 45 120 51
rect 108 39 111 45
rect 117 39 120 45
rect 108 33 120 39
rect 108 27 111 33
rect 117 27 120 33
rect 108 21 120 27
rect 108 15 111 21
rect 117 15 120 21
rect 108 9 120 15
rect 108 3 111 9
rect 117 3 120 9
rect 108 -3 120 3
rect 108 -9 111 -3
rect 117 -9 120 -3
rect 108 -15 120 -9
rect 108 -21 111 -15
rect 117 -21 120 -15
rect -60 -33 -57 -27
rect -51 -33 -48 -27
rect -60 -36 -48 -33
rect 108 -27 120 -21
rect 132 93 264 96
rect 132 87 135 93
rect 141 87 147 93
rect 153 87 159 93
rect 165 87 171 93
rect 177 87 183 93
rect 189 87 195 93
rect 201 87 207 93
rect 213 87 219 93
rect 225 87 231 93
rect 237 87 243 93
rect 249 87 255 93
rect 261 87 264 93
rect 132 84 264 87
rect 132 81 144 84
rect 132 75 135 81
rect 141 75 144 81
rect 132 69 144 75
rect 252 81 264 84
rect 252 75 255 81
rect 261 75 264 81
rect 132 63 135 69
rect 141 63 144 69
rect 132 57 144 63
rect 168 69 228 72
rect 168 63 171 69
rect 177 63 183 69
rect 189 63 195 69
rect 201 63 207 69
rect 213 63 219 69
rect 225 63 228 69
rect 168 60 228 63
rect 252 69 264 75
rect 252 63 255 69
rect 261 63 264 69
rect 132 51 135 57
rect 141 51 144 57
rect 132 45 144 51
rect 252 57 264 63
rect 252 51 255 57
rect 261 51 264 57
rect 132 39 135 45
rect 141 39 144 45
rect 132 33 144 39
rect 132 27 135 33
rect 141 27 144 33
rect 132 21 144 27
rect 132 15 135 21
rect 141 15 144 21
rect 132 9 144 15
rect 132 3 135 9
rect 141 3 144 9
rect 132 -3 144 3
rect 132 -9 135 -3
rect 141 -9 144 -3
rect 132 -12 144 -9
rect 156 45 168 48
rect 156 39 159 45
rect 165 39 168 45
rect 156 33 168 39
rect 156 27 159 33
rect 165 27 168 33
rect 156 21 168 27
rect 156 15 159 21
rect 165 15 168 21
rect 156 -12 168 15
rect 228 45 240 48
rect 228 39 231 45
rect 237 39 240 45
rect 228 33 240 39
rect 228 27 231 33
rect 237 27 240 33
rect 228 21 240 27
rect 228 15 231 21
rect 237 15 240 21
rect 228 12 240 15
rect 252 45 264 51
rect 252 39 255 45
rect 261 39 264 45
rect 252 33 264 39
rect 252 27 255 33
rect 261 27 264 33
rect 252 21 264 27
rect 252 15 255 21
rect 261 15 264 21
rect 252 9 264 15
rect 252 3 255 9
rect 261 3 264 9
rect 252 -3 264 3
rect 252 -9 255 -3
rect 261 -9 264 -3
rect 252 -12 264 -9
rect 132 -15 264 -12
rect 132 -21 135 -15
rect 141 -21 147 -15
rect 153 -21 159 -15
rect 165 -21 171 -15
rect 177 -21 183 -15
rect 189 -21 195 -15
rect 201 -21 207 -15
rect 213 -21 219 -15
rect 225 -21 231 -15
rect 237 -21 243 -15
rect 249 -21 255 -15
rect 261 -21 264 -15
rect 132 -24 264 -21
rect 276 93 288 99
rect 276 87 279 93
rect 285 87 288 93
rect 276 81 288 87
rect 276 75 279 81
rect 285 75 288 81
rect 276 69 288 75
rect 276 63 279 69
rect 285 63 288 69
rect 276 57 288 63
rect 276 51 279 57
rect 285 51 288 57
rect 276 45 288 51
rect 276 39 279 45
rect 285 39 288 45
rect 276 33 288 39
rect 276 27 279 33
rect 285 27 288 33
rect 276 21 288 27
rect 276 15 279 21
rect 285 15 288 21
rect 276 9 288 15
rect 276 3 279 9
rect 285 3 288 9
rect 276 -3 288 3
rect 276 -9 279 -3
rect 285 -9 288 -3
rect 276 -15 288 -9
rect 276 -21 279 -15
rect 285 -21 288 -15
rect 108 -33 111 -27
rect 117 -33 120 -27
rect 108 -36 120 -33
rect 276 -27 288 -21
rect 276 -33 279 -27
rect 285 -33 288 -27
rect 276 -36 288 -33
rect -60 -39 288 -36
rect -60 -45 -57 -39
rect -51 -45 -45 -39
rect -39 -45 -33 -39
rect -27 -45 -21 -39
rect -15 -45 -9 -39
rect -3 -45 3 -39
rect 9 -45 15 -39
rect 21 -45 27 -39
rect 33 -45 39 -39
rect 45 -45 51 -39
rect 57 -45 63 -39
rect 69 -45 75 -39
rect 81 -45 87 -39
rect 93 -45 99 -39
rect 105 -45 111 -39
rect 117 -45 123 -39
rect 129 -45 135 -39
rect 141 -45 147 -39
rect 153 -45 159 -39
rect 165 -45 171 -39
rect 177 -45 183 -39
rect 189 -45 195 -39
rect 201 -45 207 -39
rect 213 -45 219 -39
rect 225 -45 231 -39
rect 237 -45 243 -39
rect 249 -45 255 -39
rect 261 -45 267 -39
rect 273 -45 279 -39
rect 285 -45 288 -39
rect -60 -48 288 -45
rect -60 -51 -48 -48
rect -60 -57 -57 -51
rect -51 -57 -48 -51
rect -60 -63 -48 -57
rect 108 -51 120 -48
rect 108 -57 111 -51
rect 117 -57 120 -51
rect -60 -69 -57 -63
rect -51 -69 -48 -63
rect -60 -75 -48 -69
rect -60 -81 -57 -75
rect -51 -81 -48 -75
rect -60 -87 -48 -81
rect -60 -93 -57 -87
rect -51 -93 -48 -87
rect -60 -99 -48 -93
rect -60 -105 -57 -99
rect -51 -105 -48 -99
rect -60 -111 -48 -105
rect -60 -117 -57 -111
rect -51 -117 -48 -111
rect -60 -123 -48 -117
rect -60 -129 -57 -123
rect -51 -129 -48 -123
rect -60 -135 -48 -129
rect -60 -141 -57 -135
rect -51 -141 -48 -135
rect -60 -147 -48 -141
rect -60 -153 -57 -147
rect -51 -153 -48 -147
rect -60 -159 -48 -153
rect -60 -165 -57 -159
rect -51 -165 -48 -159
rect -60 -171 -48 -165
rect -60 -177 -57 -171
rect -51 -177 -48 -171
rect -60 -183 -48 -177
rect -36 -63 96 -60
rect -36 -69 -33 -63
rect -27 -69 -21 -63
rect -15 -69 -9 -63
rect -3 -69 3 -63
rect 9 -69 15 -63
rect 21 -69 27 -63
rect 33 -69 39 -63
rect 45 -69 51 -63
rect 57 -69 63 -63
rect 69 -69 75 -63
rect 81 -69 87 -63
rect 93 -69 96 -63
rect -36 -72 96 -69
rect -36 -75 -24 -72
rect -36 -81 -33 -75
rect -27 -81 -24 -75
rect -36 -87 -24 -81
rect -36 -93 -33 -87
rect -27 -93 -24 -87
rect -36 -99 -24 -93
rect -36 -105 -33 -99
rect -27 -105 -24 -99
rect -36 -111 -24 -105
rect -36 -117 -33 -111
rect -27 -117 -24 -111
rect -36 -123 -24 -117
rect -36 -129 -33 -123
rect -27 -129 -24 -123
rect -36 -135 -24 -129
rect -12 -99 0 -96
rect -12 -105 -9 -99
rect -3 -105 0 -99
rect -12 -111 0 -105
rect -12 -117 -9 -111
rect -3 -117 0 -111
rect -12 -123 0 -117
rect -12 -129 -9 -123
rect -3 -129 0 -123
rect -12 -132 0 -129
rect 60 -99 72 -72
rect 60 -105 63 -99
rect 69 -105 72 -99
rect 60 -111 72 -105
rect 60 -117 63 -111
rect 69 -117 72 -111
rect 60 -123 72 -117
rect 60 -129 63 -123
rect 69 -129 72 -123
rect 60 -132 72 -129
rect 84 -75 96 -72
rect 84 -81 87 -75
rect 93 -81 96 -75
rect 84 -87 96 -81
rect 84 -93 87 -87
rect 93 -93 96 -87
rect 84 -99 96 -93
rect 84 -105 87 -99
rect 93 -105 96 -99
rect 84 -111 96 -105
rect 84 -117 87 -111
rect 93 -117 96 -111
rect 84 -123 96 -117
rect 84 -129 87 -123
rect 93 -129 96 -123
rect -36 -141 -33 -135
rect -27 -141 -24 -135
rect -36 -147 -24 -141
rect 84 -135 96 -129
rect 84 -141 87 -135
rect 93 -141 96 -135
rect -36 -153 -33 -147
rect -27 -153 -24 -147
rect -36 -159 -24 -153
rect 0 -147 60 -144
rect 0 -153 3 -147
rect 9 -153 15 -147
rect 21 -153 27 -147
rect 33 -153 39 -147
rect 45 -153 51 -147
rect 57 -153 60 -147
rect 0 -156 60 -153
rect 84 -147 96 -141
rect 84 -153 87 -147
rect 93 -153 96 -147
rect -36 -165 -33 -159
rect -27 -165 -24 -159
rect -36 -168 -24 -165
rect 84 -159 96 -153
rect 84 -165 87 -159
rect 93 -165 96 -159
rect 84 -168 96 -165
rect -36 -171 96 -168
rect -36 -177 -33 -171
rect -27 -177 -21 -171
rect -15 -177 -9 -171
rect -3 -177 3 -171
rect 9 -177 15 -171
rect 21 -177 27 -171
rect 33 -177 39 -171
rect 45 -177 51 -171
rect 57 -177 63 -171
rect 69 -177 75 -171
rect 81 -177 87 -171
rect 93 -177 96 -171
rect -36 -180 96 -177
rect 108 -63 120 -57
rect 276 -51 288 -48
rect 276 -57 279 -51
rect 285 -57 288 -51
rect 108 -69 111 -63
rect 117 -69 120 -63
rect 108 -75 120 -69
rect 108 -81 111 -75
rect 117 -81 120 -75
rect 108 -87 120 -81
rect 108 -93 111 -87
rect 117 -93 120 -87
rect 108 -99 120 -93
rect 108 -105 111 -99
rect 117 -105 120 -99
rect 108 -111 120 -105
rect 108 -117 111 -111
rect 117 -117 120 -111
rect 108 -123 120 -117
rect 108 -129 111 -123
rect 117 -129 120 -123
rect 108 -135 120 -129
rect 108 -141 111 -135
rect 117 -141 120 -135
rect 108 -147 120 -141
rect 108 -153 111 -147
rect 117 -153 120 -147
rect 108 -159 120 -153
rect 108 -165 111 -159
rect 117 -165 120 -159
rect 108 -171 120 -165
rect 108 -177 111 -171
rect 117 -177 120 -171
rect -60 -189 -57 -183
rect -51 -189 -48 -183
rect -60 -192 -48 -189
rect 108 -183 120 -177
rect 132 -63 264 -60
rect 132 -69 135 -63
rect 141 -69 147 -63
rect 153 -69 159 -63
rect 165 -69 171 -63
rect 177 -69 183 -63
rect 189 -69 195 -63
rect 201 -69 207 -63
rect 213 -69 219 -63
rect 225 -69 231 -63
rect 237 -69 243 -63
rect 249 -69 255 -63
rect 261 -69 264 -63
rect 132 -72 264 -69
rect 132 -75 144 -72
rect 132 -81 135 -75
rect 141 -81 144 -75
rect 132 -87 144 -81
rect 132 -93 135 -87
rect 141 -93 144 -87
rect 132 -99 144 -93
rect 132 -105 135 -99
rect 141 -105 144 -99
rect 132 -111 144 -105
rect 132 -117 135 -111
rect 141 -117 144 -111
rect 132 -123 144 -117
rect 132 -129 135 -123
rect 141 -129 144 -123
rect 132 -135 144 -129
rect 156 -99 168 -72
rect 252 -75 264 -72
rect 252 -81 255 -75
rect 261 -81 264 -75
rect 252 -87 264 -81
rect 252 -93 255 -87
rect 261 -93 264 -87
rect 156 -105 159 -99
rect 165 -105 168 -99
rect 156 -111 168 -105
rect 156 -117 159 -111
rect 165 -117 168 -111
rect 156 -123 168 -117
rect 156 -129 159 -123
rect 165 -129 168 -123
rect 156 -132 168 -129
rect 228 -99 240 -96
rect 228 -105 231 -99
rect 237 -105 240 -99
rect 228 -111 240 -105
rect 228 -117 231 -111
rect 237 -117 240 -111
rect 228 -123 240 -117
rect 228 -129 231 -123
rect 237 -129 240 -123
rect 132 -141 135 -135
rect 141 -141 144 -135
rect 132 -147 144 -141
rect 228 -135 240 -129
rect 228 -141 231 -135
rect 237 -141 240 -135
rect 228 -144 240 -141
rect 132 -153 135 -147
rect 141 -153 144 -147
rect 132 -159 144 -153
rect 168 -147 240 -144
rect 168 -153 171 -147
rect 177 -153 183 -147
rect 189 -153 195 -147
rect 201 -153 207 -147
rect 213 -153 219 -147
rect 225 -153 231 -147
rect 237 -153 240 -147
rect 168 -156 240 -153
rect 252 -99 264 -93
rect 252 -105 255 -99
rect 261 -105 264 -99
rect 252 -111 264 -105
rect 252 -117 255 -111
rect 261 -117 264 -111
rect 252 -123 264 -117
rect 252 -129 255 -123
rect 261 -129 264 -123
rect 252 -135 264 -129
rect 252 -141 255 -135
rect 261 -141 264 -135
rect 252 -147 264 -141
rect 252 -153 255 -147
rect 261 -153 264 -147
rect 132 -165 135 -159
rect 141 -165 144 -159
rect 132 -168 144 -165
rect 252 -159 264 -153
rect 252 -165 255 -159
rect 261 -165 264 -159
rect 252 -168 264 -165
rect 132 -171 264 -168
rect 132 -177 135 -171
rect 141 -177 147 -171
rect 153 -177 159 -171
rect 165 -177 171 -171
rect 177 -177 183 -171
rect 189 -177 195 -171
rect 201 -177 207 -171
rect 213 -177 219 -171
rect 225 -177 231 -171
rect 237 -177 243 -171
rect 249 -177 255 -171
rect 261 -177 264 -171
rect 132 -180 264 -177
rect 276 -63 288 -57
rect 276 -69 279 -63
rect 285 -69 288 -63
rect 276 -75 288 -69
rect 276 -81 279 -75
rect 285 -81 288 -75
rect 276 -87 288 -81
rect 276 -93 279 -87
rect 285 -93 288 -87
rect 276 -99 288 -93
rect 276 -105 279 -99
rect 285 -105 288 -99
rect 276 -111 288 -105
rect 276 -117 279 -111
rect 285 -117 288 -111
rect 276 -123 288 -117
rect 276 -129 279 -123
rect 285 -129 288 -123
rect 276 -135 288 -129
rect 276 -141 279 -135
rect 285 -141 288 -135
rect 276 -147 288 -141
rect 276 -153 279 -147
rect 285 -153 288 -147
rect 276 -159 288 -153
rect 276 -165 279 -159
rect 285 -165 288 -159
rect 276 -171 288 -165
rect 276 -177 279 -171
rect 285 -177 288 -171
rect 108 -189 111 -183
rect 117 -189 120 -183
rect 108 -192 120 -189
rect 276 -183 288 -177
rect 276 -189 279 -183
rect 285 -189 288 -183
rect 276 -192 288 -189
rect -60 -195 288 -192
rect -60 -201 -57 -195
rect -51 -201 -45 -195
rect -39 -201 -33 -195
rect -27 -201 -21 -195
rect -15 -201 -9 -195
rect -3 -201 3 -195
rect 9 -201 15 -195
rect 21 -201 27 -195
rect 33 -201 39 -195
rect 45 -201 51 -195
rect 57 -201 63 -195
rect 69 -201 75 -195
rect 81 -201 87 -195
rect 93 -201 99 -195
rect 105 -201 111 -195
rect 117 -201 123 -195
rect 129 -201 135 -195
rect 141 -201 147 -195
rect 153 -201 159 -195
rect 165 -201 171 -195
rect 177 -201 183 -195
rect 189 -201 195 -195
rect 201 -201 207 -195
rect 213 -201 219 -195
rect 225 -201 231 -195
rect 237 -201 243 -195
rect 249 -201 255 -195
rect 261 -201 267 -195
rect 273 -201 279 -195
rect 285 -201 288 -195
rect -60 -204 288 -201
rect -60 -207 -48 -204
rect -60 -213 -57 -207
rect -51 -213 -48 -207
rect -60 -219 -48 -213
rect 108 -207 120 -204
rect 108 -213 111 -207
rect 117 -213 120 -207
rect -60 -225 -57 -219
rect -51 -225 -48 -219
rect -60 -231 -48 -225
rect -60 -237 -57 -231
rect -51 -237 -48 -231
rect -60 -243 -48 -237
rect -60 -249 -57 -243
rect -51 -249 -48 -243
rect -60 -255 -48 -249
rect -60 -261 -57 -255
rect -51 -261 -48 -255
rect -60 -267 -48 -261
rect -60 -273 -57 -267
rect -51 -273 -48 -267
rect -60 -279 -48 -273
rect -60 -285 -57 -279
rect -51 -285 -48 -279
rect -60 -291 -48 -285
rect -60 -297 -57 -291
rect -51 -297 -48 -291
rect -60 -303 -48 -297
rect -60 -309 -57 -303
rect -51 -309 -48 -303
rect -60 -315 -48 -309
rect -60 -321 -57 -315
rect -51 -321 -48 -315
rect -60 -327 -48 -321
rect -60 -333 -57 -327
rect -51 -333 -48 -327
rect -60 -339 -48 -333
rect -36 -219 96 -216
rect -36 -225 -33 -219
rect -27 -225 -21 -219
rect -15 -225 -9 -219
rect -3 -225 3 -219
rect 9 -225 15 -219
rect 21 -225 27 -219
rect 33 -225 39 -219
rect 45 -225 51 -219
rect 57 -225 63 -219
rect 69 -225 75 -219
rect 81 -225 87 -219
rect 93 -225 96 -219
rect -36 -228 96 -225
rect -36 -231 -24 -228
rect -36 -237 -33 -231
rect -27 -237 -24 -231
rect -36 -243 -24 -237
rect 84 -231 96 -228
rect 84 -237 87 -231
rect 93 -237 96 -231
rect -36 -249 -33 -243
rect -27 -249 -24 -243
rect -36 -255 -24 -249
rect -36 -261 -33 -255
rect -27 -261 -24 -255
rect -36 -267 -24 -261
rect -36 -273 -33 -267
rect -27 -273 -24 -267
rect -36 -279 -24 -273
rect -36 -285 -33 -279
rect -27 -285 -24 -279
rect -36 -291 -24 -285
rect -36 -297 -33 -291
rect -27 -297 -24 -291
rect -36 -303 -24 -297
rect -12 -243 60 -240
rect -12 -249 3 -243
rect 9 -249 15 -243
rect 21 -249 27 -243
rect 33 -249 39 -243
rect 45 -249 51 -243
rect 57 -249 60 -243
rect -12 -252 60 -249
rect 84 -243 96 -237
rect 84 -249 87 -243
rect 93 -249 96 -243
rect -12 -267 0 -252
rect 84 -255 96 -249
rect 84 -261 87 -255
rect 93 -261 96 -255
rect -12 -273 -9 -267
rect -3 -273 0 -267
rect -12 -279 0 -273
rect -12 -285 -9 -279
rect -3 -285 0 -279
rect -12 -291 0 -285
rect -12 -297 -9 -291
rect -3 -297 0 -291
rect -12 -300 0 -297
rect 60 -267 72 -264
rect 60 -273 63 -267
rect 69 -273 72 -267
rect 60 -279 72 -273
rect 60 -285 63 -279
rect 69 -285 72 -279
rect 60 -291 72 -285
rect 60 -297 63 -291
rect 69 -297 72 -291
rect -36 -309 -33 -303
rect -27 -309 -24 -303
rect -36 -315 -24 -309
rect -36 -321 -33 -315
rect -27 -321 -24 -315
rect -36 -324 -24 -321
rect 60 -324 72 -297
rect 84 -267 96 -261
rect 84 -273 87 -267
rect 93 -273 96 -267
rect 84 -279 96 -273
rect 84 -285 87 -279
rect 93 -285 96 -279
rect 84 -291 96 -285
rect 84 -297 87 -291
rect 93 -297 96 -291
rect 84 -303 96 -297
rect 84 -309 87 -303
rect 93 -309 96 -303
rect 84 -315 96 -309
rect 84 -321 87 -315
rect 93 -321 96 -315
rect 84 -324 96 -321
rect -36 -327 96 -324
rect -36 -333 -33 -327
rect -27 -333 -21 -327
rect -15 -333 -9 -327
rect -3 -333 3 -327
rect 9 -333 15 -327
rect 21 -333 27 -327
rect 33 -333 39 -327
rect 45 -333 51 -327
rect 57 -333 63 -327
rect 69 -333 75 -327
rect 81 -333 87 -327
rect 93 -333 96 -327
rect -36 -336 96 -333
rect 108 -219 120 -213
rect 108 -225 111 -219
rect 117 -225 120 -219
rect 108 -231 120 -225
rect 108 -237 111 -231
rect 117 -237 120 -231
rect 108 -243 120 -237
rect 276 -207 288 -204
rect 276 -213 279 -207
rect 285 -213 288 -207
rect 276 -219 288 -213
rect 276 -225 279 -219
rect 285 -225 288 -219
rect 276 -231 288 -225
rect 276 -237 279 -231
rect 285 -237 288 -231
rect 108 -249 111 -243
rect 117 -249 120 -243
rect 108 -255 120 -249
rect 168 -243 228 -240
rect 168 -249 171 -243
rect 177 -249 183 -243
rect 189 -249 195 -243
rect 201 -249 207 -243
rect 213 -249 219 -243
rect 225 -249 228 -243
rect 168 -252 228 -249
rect 276 -243 288 -237
rect 276 -249 279 -243
rect 285 -249 288 -243
rect 108 -261 111 -255
rect 117 -261 120 -255
rect 108 -267 120 -261
rect 276 -255 288 -249
rect 276 -261 279 -255
rect 285 -261 288 -255
rect 108 -273 111 -267
rect 117 -273 120 -267
rect 108 -279 120 -273
rect 108 -285 111 -279
rect 117 -285 120 -279
rect 108 -291 120 -285
rect 108 -297 111 -291
rect 117 -297 120 -291
rect 108 -303 120 -297
rect 156 -267 168 -264
rect 156 -273 159 -267
rect 165 -273 168 -267
rect 156 -279 168 -273
rect 156 -285 159 -279
rect 165 -285 168 -279
rect 156 -291 168 -285
rect 156 -297 159 -291
rect 165 -297 168 -291
rect 156 -300 168 -297
rect 228 -267 240 -264
rect 228 -273 231 -267
rect 237 -273 240 -267
rect 228 -279 240 -273
rect 228 -285 231 -279
rect 237 -285 240 -279
rect 228 -291 240 -285
rect 228 -297 231 -291
rect 237 -297 240 -291
rect 108 -309 111 -303
rect 117 -309 120 -303
rect 108 -315 120 -309
rect 108 -321 111 -315
rect 117 -321 120 -315
rect 108 -327 120 -321
rect 108 -333 111 -327
rect 117 -333 120 -327
rect -60 -345 -57 -339
rect -51 -345 -48 -339
rect -60 -348 -48 -345
rect 108 -339 120 -333
rect 108 -345 111 -339
rect 117 -345 120 -339
rect 108 -348 120 -345
rect 228 -348 240 -297
rect 276 -267 288 -261
rect 276 -273 279 -267
rect 285 -273 288 -267
rect 276 -279 288 -273
rect 276 -285 279 -279
rect 285 -285 288 -279
rect 276 -291 288 -285
rect 276 -297 279 -291
rect 285 -297 288 -291
rect 276 -303 288 -297
rect 276 -309 279 -303
rect 285 -309 288 -303
rect 276 -315 288 -309
rect 276 -321 279 -315
rect 285 -321 288 -315
rect 276 -327 288 -321
rect 276 -333 279 -327
rect 285 -333 288 -327
rect 276 -339 288 -333
rect 276 -345 279 -339
rect 285 -345 288 -339
rect 276 -348 288 -345
rect -60 -351 288 -348
rect -60 -357 -57 -351
rect -51 -357 -45 -351
rect -39 -357 -33 -351
rect -27 -357 -21 -351
rect -15 -357 -9 -351
rect -3 -357 3 -351
rect 9 -357 15 -351
rect 21 -357 27 -351
rect 33 -357 39 -351
rect 45 -357 51 -351
rect 57 -357 63 -351
rect 69 -357 75 -351
rect 81 -357 87 -351
rect 93 -357 99 -351
rect 105 -357 111 -351
rect 117 -357 123 -351
rect 129 -357 135 -351
rect 141 -357 147 -351
rect 153 -357 159 -351
rect 165 -357 171 -351
rect 177 -357 183 -351
rect 189 -357 195 -351
rect 201 -357 207 -351
rect 213 -357 219 -351
rect 225 -357 231 -351
rect 237 -357 243 -351
rect 249 -357 255 -351
rect 261 -357 267 -351
rect 273 -357 279 -351
rect 285 -357 288 -351
rect -60 -360 288 -357
<< via1 >>
rect 231 111 237 117
rect -57 -21 -51 -15
rect -33 87 -27 93
rect -33 75 -27 81
rect -33 63 -27 69
rect -33 51 -27 57
rect -33 39 -27 45
rect -33 27 -27 33
rect -33 15 -27 21
rect -9 63 -3 69
rect -9 51 -3 57
rect -33 3 -27 9
rect -33 -9 -27 -3
rect -33 -21 -27 -15
rect 135 87 141 93
rect 135 75 141 81
rect 135 63 141 69
rect 195 63 201 69
rect 135 51 141 57
rect 135 39 141 45
rect 135 27 141 33
rect 135 15 141 21
rect 135 3 141 9
rect 135 -9 141 -3
rect 231 39 237 45
rect 231 27 237 33
rect 231 15 237 21
rect 135 -21 141 -15
rect 279 -21 285 -15
rect -57 -69 -51 -63
rect 87 -69 93 -63
rect -9 -105 -3 -99
rect -9 -117 -3 -111
rect -9 -129 -3 -123
rect 87 -81 93 -75
rect 87 -93 93 -87
rect 87 -105 93 -99
rect 87 -117 93 -111
rect 87 -129 93 -123
rect 87 -141 93 -135
rect 27 -153 33 -147
rect 87 -153 93 -147
rect 87 -165 93 -159
rect 87 -177 93 -171
rect 255 -69 261 -63
rect 255 -81 261 -75
rect 255 -93 261 -87
rect 231 -141 237 -135
rect 231 -153 237 -147
rect 255 -105 261 -99
rect 255 -117 261 -111
rect 255 -129 261 -123
rect 255 -141 261 -135
rect 255 -153 261 -147
rect 255 -165 261 -159
rect 255 -177 261 -171
rect 279 -69 285 -63
rect -9 -201 -3 -195
rect -57 -333 -51 -327
rect -33 -225 -27 -219
rect -33 -237 -27 -231
rect -33 -249 -27 -243
rect -33 -261 -27 -255
rect -33 -273 -27 -267
rect -33 -285 -27 -279
rect -33 -297 -27 -291
rect 3 -249 9 -243
rect 15 -249 21 -243
rect 27 -249 33 -243
rect 39 -249 45 -243
rect 51 -249 57 -243
rect -33 -309 -27 -303
rect -33 -321 -27 -315
rect -33 -333 -27 -327
rect 171 -249 177 -243
rect 183 -249 189 -243
rect 195 -249 201 -243
rect 207 -249 213 -243
rect 219 -249 225 -243
rect 159 -273 165 -267
rect 111 -333 117 -327
rect -57 -345 -51 -339
rect 111 -345 117 -339
rect 279 -333 285 -327
rect 279 -345 285 -339
rect -57 -357 -51 -351
rect 111 -357 117 -351
rect 279 -357 285 -351
<< metal2 >>
rect -36 117 -24 120
rect -36 111 -33 117
rect -27 111 -24 117
rect -36 105 -24 111
rect -36 99 -33 105
rect -27 99 -24 105
rect -36 93 -24 99
rect 228 117 240 120
rect 228 111 231 117
rect 237 111 240 117
rect -36 87 -33 93
rect -27 87 -24 93
rect -36 81 -24 87
rect -36 75 -33 81
rect -27 75 -24 81
rect -36 69 -24 75
rect 132 93 144 96
rect 132 87 135 93
rect 141 87 144 93
rect 132 81 144 87
rect 132 75 135 81
rect 141 75 144 81
rect -36 63 -33 69
rect -27 63 -24 69
rect -36 57 -24 63
rect -36 51 -33 57
rect -27 51 -24 57
rect -36 45 -24 51
rect -36 39 -33 45
rect -27 39 -24 45
rect -36 33 -24 39
rect -36 27 -33 33
rect -27 27 -24 33
rect -36 21 -24 27
rect -36 15 -33 21
rect -27 15 -24 21
rect -36 9 -24 15
rect -36 3 -33 9
rect -27 3 -24 9
rect -36 -3 -24 3
rect -36 -9 -33 -3
rect -27 -9 -24 -3
rect -60 -15 -48 -12
rect -60 -21 -57 -15
rect -51 -21 -48 -15
rect -60 -63 -48 -21
rect -60 -69 -57 -63
rect -51 -69 -48 -63
rect -60 -327 -48 -69
rect -60 -333 -57 -327
rect -51 -333 -48 -327
rect -60 -339 -48 -333
rect -36 -15 -24 -9
rect -36 -21 -33 -15
rect -27 -21 -24 -15
rect -36 -171 -24 -21
rect -12 69 0 72
rect -12 63 -9 69
rect -3 63 0 69
rect -12 57 0 63
rect -12 51 -9 57
rect -3 51 0 57
rect -12 -39 0 51
rect 108 69 120 72
rect 108 63 111 69
rect 117 63 120 69
rect -12 -45 -9 -39
rect -3 -45 0 -39
rect -12 -48 0 -45
rect 84 -39 96 -36
rect 84 -45 87 -39
rect 93 -45 96 -39
rect 84 -63 96 -45
rect 84 -69 87 -63
rect 93 -69 96 -63
rect 84 -75 96 -69
rect 84 -81 87 -75
rect 93 -81 96 -75
rect 84 -87 96 -81
rect 84 -93 87 -87
rect 93 -93 96 -87
rect -36 -177 -33 -171
rect -27 -177 -24 -171
rect -36 -183 -24 -177
rect -36 -189 -33 -183
rect -27 -189 -24 -183
rect -36 -195 -24 -189
rect -36 -201 -33 -195
rect -27 -201 -24 -195
rect -36 -219 -24 -201
rect -12 -99 0 -96
rect -12 -105 -9 -99
rect -3 -105 0 -99
rect -12 -111 0 -105
rect -12 -117 -9 -111
rect -3 -117 0 -111
rect -12 -123 0 -117
rect -12 -129 -9 -123
rect -3 -129 0 -123
rect -12 -195 0 -129
rect 84 -99 96 -93
rect 84 -105 87 -99
rect 93 -105 96 -99
rect 84 -111 96 -105
rect 84 -117 87 -111
rect 93 -117 96 -111
rect 84 -123 96 -117
rect 84 -129 87 -123
rect 93 -129 96 -123
rect 84 -135 96 -129
rect 84 -141 87 -135
rect 93 -141 96 -135
rect 24 -147 36 -144
rect 24 -153 27 -147
rect 33 -153 36 -147
rect 24 -156 36 -153
rect 84 -147 96 -141
rect 84 -153 87 -147
rect 93 -153 96 -147
rect 84 -159 96 -153
rect 84 -165 87 -159
rect 93 -165 96 -159
rect 84 -171 96 -165
rect 84 -177 87 -171
rect 93 -177 96 -171
rect 84 -180 96 -177
rect 108 -147 120 63
rect 132 69 144 75
rect 132 63 135 69
rect 141 63 144 69
rect 132 57 144 63
rect 192 69 204 72
rect 192 63 195 69
rect 201 63 204 69
rect 192 60 204 63
rect 132 51 135 57
rect 141 51 144 57
rect 132 45 144 51
rect 132 39 135 45
rect 141 39 144 45
rect 132 33 144 39
rect 132 27 135 33
rect 141 27 144 33
rect 132 21 144 27
rect 132 15 135 21
rect 141 15 144 21
rect 132 9 144 15
rect 228 45 240 111
rect 228 39 231 45
rect 237 39 240 45
rect 228 33 240 39
rect 228 27 231 33
rect 237 27 240 33
rect 228 21 240 27
rect 228 15 231 21
rect 237 15 240 21
rect 228 12 240 15
rect 252 117 264 120
rect 252 111 255 117
rect 261 111 264 117
rect 252 105 264 111
rect 252 99 255 105
rect 261 99 264 105
rect 252 93 264 99
rect 252 87 255 93
rect 261 87 264 93
rect 132 3 135 9
rect 141 3 144 9
rect 132 -3 144 3
rect 132 -9 135 -3
rect 141 -9 144 -3
rect 132 -15 144 -9
rect 132 -21 135 -15
rect 141 -21 144 -15
rect 132 -39 144 -21
rect 132 -45 135 -39
rect 141 -45 144 -39
rect 132 -48 144 -45
rect 228 -39 240 -36
rect 228 -45 231 -39
rect 237 -45 240 -39
rect 108 -153 111 -147
rect 117 -153 120 -147
rect -12 -201 -9 -195
rect -3 -201 0 -195
rect -12 -204 0 -201
rect -36 -225 -33 -219
rect -27 -225 -24 -219
rect -36 -231 -24 -225
rect -36 -237 -33 -231
rect -27 -237 -24 -231
rect -36 -243 -24 -237
rect -36 -249 -33 -243
rect -27 -249 -24 -243
rect -36 -255 -24 -249
rect 0 -243 60 -240
rect 0 -249 3 -243
rect 9 -249 15 -243
rect 21 -249 27 -243
rect 33 -249 39 -243
rect 45 -249 51 -243
rect 57 -249 60 -243
rect 0 -252 60 -249
rect -36 -261 -33 -255
rect -27 -261 -24 -255
rect -36 -267 -24 -261
rect -36 -273 -33 -267
rect -27 -273 -24 -267
rect -36 -279 -24 -273
rect 108 -267 120 -153
rect 228 -135 240 -45
rect 228 -141 231 -135
rect 237 -141 240 -135
rect 228 -147 240 -141
rect 228 -153 231 -147
rect 237 -153 240 -147
rect 228 -156 240 -153
rect 252 -63 264 87
rect 252 -69 255 -63
rect 261 -69 264 -63
rect 252 -75 264 -69
rect 252 -81 255 -75
rect 261 -81 264 -75
rect 252 -87 264 -81
rect 252 -93 255 -87
rect 261 -93 264 -87
rect 252 -99 264 -93
rect 252 -105 255 -99
rect 261 -105 264 -99
rect 252 -111 264 -105
rect 252 -117 255 -111
rect 261 -117 264 -111
rect 252 -123 264 -117
rect 252 -129 255 -123
rect 261 -129 264 -123
rect 252 -135 264 -129
rect 252 -141 255 -135
rect 261 -141 264 -135
rect 252 -147 264 -141
rect 252 -153 255 -147
rect 261 -153 264 -147
rect 252 -159 264 -153
rect 252 -165 255 -159
rect 261 -165 264 -159
rect 252 -171 264 -165
rect 252 -177 255 -171
rect 261 -177 264 -171
rect 252 -183 264 -177
rect 252 -189 255 -183
rect 261 -189 264 -183
rect 132 -204 144 -192
rect 252 -195 264 -189
rect 252 -201 255 -195
rect 261 -201 264 -195
rect 252 -204 264 -201
rect 276 -15 288 -12
rect 276 -21 279 -15
rect 285 -21 288 -15
rect 276 -63 288 -21
rect 276 -69 279 -63
rect 285 -69 288 -63
rect 168 -243 228 -240
rect 168 -249 171 -243
rect 177 -249 183 -243
rect 189 -249 195 -243
rect 201 -249 207 -243
rect 213 -249 219 -243
rect 225 -249 228 -243
rect 168 -252 228 -249
rect 108 -273 111 -267
rect 117 -273 120 -267
rect 108 -276 120 -273
rect 156 -267 168 -264
rect 156 -273 159 -267
rect 165 -273 168 -267
rect 156 -276 168 -273
rect -36 -285 -33 -279
rect -27 -285 -24 -279
rect -36 -291 -24 -285
rect -36 -297 -33 -291
rect -27 -297 -24 -291
rect -36 -303 -24 -297
rect -36 -309 -33 -303
rect -27 -309 -24 -303
rect -36 -315 -24 -309
rect -36 -321 -33 -315
rect -27 -321 -24 -315
rect -36 -327 -24 -321
rect -36 -333 -33 -327
rect -27 -333 -24 -327
rect -36 -336 -24 -333
rect 108 -327 120 -324
rect 108 -333 111 -327
rect 117 -333 120 -327
rect -60 -345 -57 -339
rect -51 -345 -48 -339
rect -60 -351 -48 -345
rect -60 -357 -57 -351
rect -51 -357 -48 -351
rect -60 -360 -48 -357
rect 108 -339 120 -333
rect 108 -345 111 -339
rect 117 -345 120 -339
rect 108 -351 120 -345
rect 108 -357 111 -351
rect 117 -357 120 -351
rect 108 -360 120 -357
rect 276 -327 288 -69
rect 276 -333 279 -327
rect 285 -333 288 -327
rect 276 -339 288 -333
rect 276 -345 279 -339
rect 285 -345 288 -339
rect 276 -351 288 -345
rect 276 -357 279 -351
rect 285 -357 288 -351
rect 276 -360 288 -357
<< via2 >>
rect -33 111 -27 117
rect -33 99 -27 105
rect -33 87 -27 93
rect -57 -21 -51 -15
rect -57 -69 -51 -63
rect -57 -333 -51 -327
rect 111 63 117 69
rect -9 -45 -3 -39
rect 87 -45 93 -39
rect -33 -177 -27 -171
rect -33 -189 -27 -183
rect -33 -201 -27 -195
rect 27 -153 33 -147
rect 195 63 201 69
rect 255 111 261 117
rect 255 99 261 105
rect 255 87 261 93
rect 135 -45 141 -39
rect 231 -45 237 -39
rect 111 -153 117 -147
rect 3 -249 9 -243
rect 15 -249 21 -243
rect 27 -249 33 -243
rect 39 -249 45 -243
rect 51 -249 57 -243
rect 255 -177 261 -171
rect 255 -189 261 -183
rect 255 -201 261 -195
rect 279 -21 285 -15
rect 279 -69 285 -63
rect 171 -249 177 -243
rect 183 -249 189 -243
rect 195 -249 201 -243
rect 207 -249 213 -243
rect 219 -249 225 -243
rect 111 -273 117 -267
rect 159 -273 165 -267
rect 111 -333 117 -327
rect -57 -345 -51 -339
rect -57 -357 -51 -351
rect 111 -345 117 -339
rect 111 -357 117 -351
rect 279 -333 285 -327
rect 279 -345 285 -339
rect 279 -357 285 -351
<< metal3 >>
rect -60 117 288 120
rect -60 111 -33 117
rect -27 111 255 117
rect 261 111 288 117
rect -60 105 288 111
rect -60 99 -33 105
rect -27 99 255 105
rect 261 99 288 105
rect -60 93 288 99
rect -60 87 -33 93
rect -27 87 255 93
rect 261 87 288 93
rect -60 84 288 87
rect 108 69 228 72
rect 108 63 111 69
rect 117 63 195 69
rect 201 63 228 69
rect 108 60 228 63
rect -60 -15 288 -12
rect -60 -21 -57 -15
rect -51 -21 279 -15
rect 285 -21 288 -15
rect -60 -24 288 -21
rect -60 -39 288 -36
rect -60 -45 -9 -39
rect -3 -45 87 -39
rect 93 -45 135 -39
rect 141 -45 231 -39
rect 237 -45 288 -39
rect -60 -48 288 -45
rect -60 -63 288 -60
rect -60 -69 -57 -63
rect -51 -69 279 -63
rect 285 -69 288 -63
rect -60 -72 288 -69
rect 0 -147 120 -144
rect 0 -153 27 -147
rect 33 -153 111 -147
rect 117 -153 120 -147
rect 0 -156 120 -153
rect -60 -171 288 -168
rect -60 -177 -33 -171
rect -27 -177 255 -171
rect 261 -177 288 -171
rect -60 -183 288 -177
rect -60 -189 -33 -183
rect -27 -189 255 -183
rect 261 -189 288 -183
rect -60 -195 288 -189
rect -60 -201 -33 -195
rect -27 -201 255 -195
rect 261 -201 288 -195
rect -60 -204 288 -201
rect -12 -243 228 -240
rect -12 -249 3 -243
rect 9 -249 15 -243
rect 21 -249 27 -243
rect 33 -249 39 -243
rect 45 -249 51 -243
rect 57 -249 171 -243
rect 177 -249 183 -243
rect 189 -249 195 -243
rect 201 -249 207 -243
rect 213 -249 219 -243
rect 225 -249 228 -243
rect -12 -252 228 -249
rect 108 -267 168 -264
rect 108 -273 111 -267
rect 117 -273 159 -267
rect 165 -273 168 -267
rect 108 -276 168 -273
rect -60 -327 288 -324
rect -60 -333 -57 -327
rect -51 -333 111 -327
rect 117 -333 279 -327
rect 285 -333 288 -327
rect -60 -339 288 -333
rect -60 -345 -57 -339
rect -51 -345 111 -339
rect 117 -345 279 -339
rect 285 -345 288 -339
rect -60 -351 288 -345
rect -60 -357 -57 -351
rect -51 -357 111 -351
rect 117 -357 279 -351
rect 285 -357 288 -351
rect -60 -360 288 -357
<< labels >>
rlabel metal3 -60 -48 288 -36 0 ref
port 1 nsew
rlabel metal3 -60 84 288 120 0 vdd
port 2 nsew
rlabel metal3 -60 -360 288 -324 0 vss
port 3 nsew
rlabel metal3 132 -276 144 -264 0 tilo
rlabel metal3 132 -252 144 -240 0 tihi
<< end >>
